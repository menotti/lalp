-- IEEE Libraries -- 
library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 

entity block_ram_in is 
generic( 
        data_width : integer := 8; 
        address_width : integer := 8 
); 
port( 
        data_in : in std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        address : in std_logic_vector(address_width-1 downto 0); 
        we: in std_logic := '0'; 
        oe: in std_logic := '1'; 
        clk : in std_logic; 
        data_out : out std_logic_vector(data_width-1 downto 0)); 
end block_ram_in; 

architecture rtl of block_ram_in is 

constant mem_depth : integer := 2**address_width; 
type ram_type is array (mem_depth-1 downto 0) 
of std_logic_vector (data_width-1 downto 0); 

signal read_a : std_logic_vector(address_width-1 downto 0); 
signal RAM : ram_type := ram_type'( 
	 ("00000100000000000000000000000000"),	 -- 127	0
	 ("00000010000000000000000000000000"),	 -- 126	0
	 ("00000001000000000000000000000000"),	 -- 125	0
	 ("00000000100000000000000000000000"),	 -- 124	0
	 ("00000000010000000000000000000000"),	 -- 123	0
	 ("00000000001000000000000000000000"),	 -- 122	0
	 ("00000000000100000000000000000000"),	 -- 121	0
	 ("00000000000000000000000000000000"),	 -- 120	0
	 ("00000000000011000000000000000000"),	 -- 119	0
	 ("00000000000000000000000000000000"),	 -- 118	0
	 ("00000000000000100000000000000000"),	 -- 117	0
	 ("00000000000000010000000000000000"),	 -- 116	0
	 ("00000000000000001000000000000000"),	 -- 115	0
	 ("00000000000000000100000000000000"),	 -- 114	0
	 ("00000000000000000010000000000000"),	 -- 113	0
	 ("00000000000000000001000000000000"),	 -- 112	0
	 ("00000000000000000000100000000000"),	 -- 111	0
	 ("00000000000000000000010000000000"),	 -- 110	0
	 ("00000000000000000000001000000000"),	 -- 109	0
	 ("00000000000000000000000100000000"),	 -- 108	0
	 ("00000000000000000000000010000000"),	 -- 107	0
	 ("00000000000000000000000001000000"),	 -- 106	0
	 ("00000000000000000000000000000000"),	 -- 105	0
	 ("00000000000000000000000000000000"),	 -- 104	0
	 ("00000000000000000000000000000000"),	 -- 103	0
	 ("00000000000000000000000000000000"),	 -- 102	0
	 ("00000000000000000000000000000000"),	 -- 101	0
	 ("00000000000000000000000000000000"),	 -- 100	0
	 ("00000000000000000000000001100011"),	 -- 99	99
	 ("00000000000000000000000000100110"),	 -- 98	38
	 ("00000000000000000000000001100001"),	 -- 97	97
	 ("00000000000000000000000001100000"),	 -- 96	96
	 ("00000000000000000000000001011111"),	 -- 95	95
	 ("00000000000000000000000001011110"),	 -- 94	94
	 ("00000000000000000000000001011101"),	 -- 93	93
	 ("00000000000000000000000001011100"),	 -- 92	92
	 ("00000000000000000000000001100000"),	 -- 91	96
	 ("00000000000000000000000001011111"),	 -- 90	95
	 ("00000000000000000000000001011001"),	 -- 89	89
	 ("00000000000000000000000000011100"),	 -- 88	28
	 ("00000000000000000000000001010111"),	 -- 87	87
	 ("00000000000000000000000001010110"),	 -- 86	86
	 ("00000000000000000000000001010101"),	 -- 85	85
	 ("00000000000000000000000001010100"),	 -- 84	84
	 ("00000000000000000000000001010011"),	 -- 83	83
	 ("00000000000000000000000001010010"),	 -- 82	82
	 ("00000000000000000000000001010111"),	 -- 81	87
	 ("00000000000000000000000001010100"),	 -- 80	84
	 ("00000000000000000000000000011101"),	 -- 79	29
	 ("00000000000000000000000000010010"),	 -- 78	18
	 ("00000000000000000000000000100101"),	 -- 77	37
	 ("00000000000000000000000001100000"),	 -- 76	96
	 ("00000000000000000000000000110111"),	 -- 75	55
	 ("00000000000000000000000000100010"),	 -- 74	34
	 ("00000000000000000000000001010011"),	 -- 73	83
	 ("00000000000000000000000001001000"),	 -- 72	72
	 ("00000000000000000000000001000100"),	 -- 71	68
	 ("00000000000000000000000000110101"),	 -- 70	53
	 ("00000000000000000000000001000101"),	 -- 69	69
	 ("00000000000000000000000001000100"),	 -- 68	68
	 ("00000000000000000000000001000011"),	 -- 67	67
	 ("00000000000000000000000001000000"),	 -- 66	64
	 ("00000000000000000000000001000001"),	 -- 65	65
	 ("00000000000000000000000001000000"),	 -- 64	64
	 ("00000000000000000000000001000010"),	 -- 63	66
	 ("00000000000000000000000000111110"),	 -- 62	62
	 ("00000000000000000000000001000101"),	 -- 61	69
	 ("00000000000000000000000000111100"),	 -- 60	60
	 ("00000000000000000000000000011101"),	 -- 59	29
	 ("00000000000000000000000000010010"),	 -- 58	18
	 ("00000000000000000000000000100101"),	 -- 57	37
	 ("00000000000000000000000001100000"),	 -- 56	96
	 ("00000000000000000000000000101101"),	 -- 55	45
	 ("00000000000000000000000000100010"),	 -- 54	34
	 ("00000000000000000000000001010011"),	 -- 53	83
	 ("00000000000000000000000001010010"),	 -- 52	82
	 ("00000000000000000000000000111100"),	 -- 51	60
	 ("00000000000000000000000000110100"),	 -- 50	52
	 ("00000000000000000000000001011001"),	 -- 49	89
	 ("00000000000000000000000000110000"),	 -- 48	48
	 ("00000000000000000000000000101111"),	 -- 47	47
	 ("00000000000000000000000000101110"),	 -- 46	46
	 ("00000000000000000000000000101101"),	 -- 45	45
	 ("00000000000000000000000000101100"),	 -- 44	44
	 ("00000000000000000000000001001001"),	 -- 43	73
	 ("00000000000000000000000000101010"),	 -- 42	42
	 ("00000000000000000000000000101001"),	 -- 41	41
	 ("00000000000000000000000000101000"),	 -- 40	40
	 ("00000000000000000000000000011101"),	 -- 39	29
	 ("00000000000000000000000000010010"),	 -- 38	18
	 ("00000000000000000000000001100001"),	 -- 37	97
	 ("00000000000000000000000001100000"),	 -- 36	96
	 ("00000000000000000000000000101101"),	 -- 35	45
	 ("00000000000000000000000000100010"),	 -- 34	34
	 ("00000000000000000000000001010011"),	 -- 33	83
	 ("00000000000000000000000001001000"),	 -- 32	72
	 ("00000000000000000000000000001100"),	 -- 31	12
	 ("00000000000000000000000000110110"),	 -- 30	54
	 ("00000000000000000000000000011101"),	 -- 29	29
	 ("00000000000000000000000000011100"),	 -- 28	28
	 ("00000000000000000000000000011011"),	 -- 27	27
	 ("00000000000000000000000000011010"),	 -- 26	26
	 ("00000000000000000000000000011001"),	 -- 25	25
	 ("00000000000000000000000000010100"),	 -- 24	20
	 ("00000000000000000000000000010111"),	 -- 23	23
	 ("00000000000000000000000001010010"),	 -- 22	82
	 ("00000000000000000000000000010111"),	 -- 21	23
	 ("00000000000000000000000000010100"),	 -- 20	20
	 ("00000000000000000000000000100111"),	 -- 19	39
	 ("00000000000000000000000000010010"),	 -- 18	18
	 ("00000000000000000000000000010001"),	 -- 17	17
	 ("00000000000000000000000000010000"),	 -- 16	16
	 ("00000000000000000000000000001111"),	 -- 15	15
	 ("00000000000000000000000000001110"),	 -- 14	14
	 ("00000000000000000000000000001101"),	 -- 13	13
	 ("00000000000000000000000001001000"),	 -- 12	72
	 ("00000000000000000000000000001110"),	 -- 11	14
	 ("00000000000000000000000000001110"),	 -- 10	14
	 ("00000000000000000000000000011101"),	 -- 9	29
	 ("00000000000000000000000000010010"),	 -- 8	18
	 ("00000000000000000000000001000011"),	 -- 7	67
	 ("00000000000000000000000001100000"),	 -- 6	96
	 ("00000000000000000000000000101101"),	 -- 5	45
	 ("00000000000000000000000000100010"),	 -- 4	34
	 ("00000000000000000000000001010011"),	 -- 3	83
	 ("00000000000000000000000000111110"),	 -- 2	62
	 ("00000000000000000000000001000001"),	 -- 1	65
	 ("00000000000000000000000000110010"));	 -- 0	50


begin 
       process (clk) 
       begin 
              if (clk'event and clk = '1') then 
                  if (we = '1') then 
                        RAM(conv_integer(address)) <= data_in; 
                        data_out <= RAM(conv_integer(read_a)); 
                  elsif (oe = '1') then 
                        data_out <= RAM(conv_integer(read_a)); 
                  end if; 
                  read_a <= address; 
             end if; 
       end process; 
end rtl; 

