library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 
entity dotprod is 
   port ( 
           \clear\  : in	 std_logic; 
           \clk\    : in	 std_logic; 
           \done\   : out std_logic; 
           \init\   : in	 std_logic; 
           \reset\  : in	 std_logic; 
           \result\ : out std_logic_vector(31 downto 0) 
); 
end dotprod; 

architecture behavior of dotprod is 

component add_op_s 
generic ( 
        w_in1	: integer := 8; 
        w_in2	: integer := 8; 
        w_out	: integer := 16 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component add_reg_op_s 
generic ( 
        w_in1	: integer := 16; 
        w_in2	: integer := 16; 
        w_out	: integer := 32; 
        initial	: integer := 0
); 
port ( 
        clk         : in	std_logic; 
        reset       : in	std_logic; 
        we          : in	std_logic := '1'; 
        Sel1        : in	std_logic_vector(0 downto 0) := "1"; 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component block_ram_a 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_107 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_115 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_123 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_131 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_139 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_147 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_155 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_163 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_171 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_179 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_187 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_19 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_195 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_203 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_211 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_219 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_227 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_235 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_243 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_251 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_259 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_27 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_35 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_43 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_51 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_59 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_67 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_75 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_83 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_91 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_a_99 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_100 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_108 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_116 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_124 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_132 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_140 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_148 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_156 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_164 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_172 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_180 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_188 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_196 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_20 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_204 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_212 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_220 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_228 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_236 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_244 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_252 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_260 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_28 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_36 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_44 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_52 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_60 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_68 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_76 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_84 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_b_92 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component counter 
generic (
        bits		: integer := 8;
        steps		: integer := 1;
        increment           : integer := 1;
        down                : integer := 0;
        condition           : integer := 0
);
port (
        input		: in	std_logic_vector(bits-1 downto 0);
        termination         : in	std_logic_vector(bits-1 downto 0);
        clk                 : in	std_logic;
        clk_en		: in	std_logic := '1';
        reset		: in	std_logic;
        load		: in	std_logic := '0';
        step		: out	std_logic;
        done		: out	std_logic;
        output		: out	std_logic_vector(bits-1 downto 0)
); 
end component; 

component delay_op 
generic ( 
        bits        : integer := 8; 
        delay       : integer := 1 
); 
port ( 
        a		: in	std_logic_vector(bits-1 downto 0); 
        clk		: in	std_logic; 
        reset	: in	std_logic; 
        a_delayed	: out	std_logic_vector(bits-1 downto 0) := (others=>'0') 
); 
end component; 

component mult_op_s 
generic ( 
        w_in1	: integer := 8; 
        w_in2	: integer := 8; 
        w_out	: integer := 16 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component reg_op 
generic ( 
        w_in	: integer := 16; 
        initial	: integer := 0 
); 
port ( 
        clk         : in	std_logic; 
        reset       : in	std_logic; 
        we          : in	std_logic := '1'; 
        I0          : in	std_logic_vector(w_in-1 downto 0); 
        O0          : out	std_logic_vector(w_in-1 downto 0) 
); 
end component; 

signal s216	: std_logic_vector(31 downto 0); 
signal s1	: std_logic_vector(31 downto 0); 
signal s352	: std_logic_vector(31 downto 0); 
signal s3	: std_logic_vector(31 downto 0); 
signal s4	: std_logic_vector(31 downto 0); 
signal s5	: std_logic_vector(31 downto 0); 
signal s7	: std_logic_vector(31 downto 0); 
signal s8	: std_logic_vector(31 downto 0); 
signal s353	: std_logic_vector(31 downto 0); 
signal s10	: std_logic_vector(31 downto 0); 
signal s11	: std_logic_vector(31 downto 0); 
signal s12	: std_logic_vector(31 downto 0); 
signal s14	: std_logic_vector(31 downto 0); 
signal s15	: std_logic_vector(31 downto 0); 
signal s354	: std_logic_vector(31 downto 0); 
signal s17	: std_logic_vector(31 downto 0); 
signal s18	: std_logic_vector(31 downto 0); 
signal s19	: std_logic_vector(31 downto 0); 
signal s21	: std_logic_vector(31 downto 0); 
signal s22	: std_logic_vector(31 downto 0); 
signal s355	: std_logic_vector(31 downto 0); 
signal s24	: std_logic_vector(31 downto 0); 
signal s25	: std_logic_vector(31 downto 0); 
signal s26	: std_logic_vector(31 downto 0); 
signal s28	: std_logic_vector(31 downto 0); 
signal s29	: std_logic_vector(31 downto 0); 
signal s356	: std_logic_vector(31 downto 0); 
signal s31	: std_logic_vector(31 downto 0); 
signal s32	: std_logic_vector(31 downto 0); 
signal s33	: std_logic_vector(31 downto 0); 
signal s35	: std_logic_vector(31 downto 0); 
signal s36	: std_logic_vector(31 downto 0); 
signal s357	: std_logic_vector(31 downto 0); 
signal s38	: std_logic_vector(31 downto 0); 
signal s39	: std_logic_vector(31 downto 0); 
signal s40	: std_logic_vector(31 downto 0); 
signal s42	: std_logic_vector(31 downto 0); 
signal s43	: std_logic_vector(31 downto 0); 
signal s358	: std_logic_vector(31 downto 0); 
signal s45	: std_logic_vector(31 downto 0); 
signal s46	: std_logic_vector(31 downto 0); 
signal s47	: std_logic_vector(31 downto 0); 
signal s49	: std_logic_vector(31 downto 0); 
signal s50	: std_logic_vector(31 downto 0); 
signal s359	: std_logic_vector(31 downto 0); 
signal s52	: std_logic_vector(31 downto 0); 
signal s53	: std_logic_vector(31 downto 0); 
signal s54	: std_logic_vector(31 downto 0); 
signal s56	: std_logic_vector(31 downto 0); 
signal s57	: std_logic_vector(31 downto 0); 
signal s360	: std_logic_vector(31 downto 0); 
signal s59	: std_logic_vector(31 downto 0); 
signal s60	: std_logic_vector(31 downto 0); 
signal s61	: std_logic_vector(31 downto 0); 
signal s63	: std_logic_vector(31 downto 0); 
signal s64	: std_logic_vector(31 downto 0); 
signal s361	: std_logic_vector(31 downto 0); 
signal s66	: std_logic_vector(31 downto 0); 
signal s67	: std_logic_vector(31 downto 0); 
signal s68	: std_logic_vector(31 downto 0); 
signal s70	: std_logic_vector(31 downto 0); 
signal s71	: std_logic_vector(31 downto 0); 
signal s362	: std_logic_vector(31 downto 0); 
signal s73	: std_logic_vector(31 downto 0); 
signal s74	: std_logic_vector(31 downto 0); 
signal s75	: std_logic_vector(31 downto 0); 
signal s77	: std_logic_vector(31 downto 0); 
signal s78	: std_logic_vector(31 downto 0); 
signal s363	: std_logic_vector(31 downto 0); 
signal s80	: std_logic_vector(31 downto 0); 
signal s81	: std_logic_vector(31 downto 0); 
signal s82	: std_logic_vector(31 downto 0); 
signal s84	: std_logic_vector(31 downto 0); 
signal s85	: std_logic_vector(31 downto 0); 
signal s364	: std_logic_vector(31 downto 0); 
signal s87	: std_logic_vector(31 downto 0); 
signal s88	: std_logic_vector(31 downto 0); 
signal s89	: std_logic_vector(31 downto 0); 
signal s91	: std_logic_vector(31 downto 0); 
signal s92	: std_logic_vector(31 downto 0); 
signal s365	: std_logic_vector(31 downto 0); 
signal s94	: std_logic_vector(31 downto 0); 
signal s95	: std_logic_vector(31 downto 0); 
signal s96	: std_logic_vector(31 downto 0); 
signal s98	: std_logic_vector(31 downto 0); 
signal s99	: std_logic_vector(31 downto 0); 
signal s366	: std_logic_vector(31 downto 0); 
signal s101	: std_logic_vector(31 downto 0); 
signal s102	: std_logic_vector(31 downto 0); 
signal s103	: std_logic_vector(31 downto 0); 
signal s105	: std_logic_vector(31 downto 0); 
signal s106	: std_logic_vector(31 downto 0); 
signal s367	: std_logic_vector(31 downto 0); 
signal s108	: std_logic_vector(31 downto 0); 
signal s109	: std_logic_vector(31 downto 0); 
signal s110	: std_logic_vector(31 downto 0); 
signal s112	: std_logic_vector(31 downto 0); 
signal s113	: std_logic_vector(31 downto 0); 
signal s368	: std_logic_vector(31 downto 0); 
signal s115	: std_logic_vector(31 downto 0); 
signal s116	: std_logic_vector(31 downto 0); 
signal s117	: std_logic_vector(31 downto 0); 
signal s119	: std_logic_vector(31 downto 0); 
signal s120	: std_logic_vector(31 downto 0); 
signal s369	: std_logic_vector(31 downto 0); 
signal s122	: std_logic_vector(31 downto 0); 
signal s123	: std_logic_vector(31 downto 0); 
signal s124	: std_logic_vector(31 downto 0); 
signal s126	: std_logic_vector(31 downto 0); 
signal s127	: std_logic_vector(31 downto 0); 
signal s370	: std_logic_vector(31 downto 0); 
signal s129	: std_logic_vector(31 downto 0); 
signal s130	: std_logic_vector(31 downto 0); 
signal s131	: std_logic_vector(31 downto 0); 
signal s133	: std_logic_vector(31 downto 0); 
signal s134	: std_logic_vector(31 downto 0); 
signal s371	: std_logic_vector(31 downto 0); 
signal s136	: std_logic_vector(31 downto 0); 
signal s137	: std_logic_vector(31 downto 0); 
signal s138	: std_logic_vector(31 downto 0); 
signal s140	: std_logic_vector(31 downto 0); 
signal s141	: std_logic_vector(31 downto 0); 
signal s372	: std_logic_vector(31 downto 0); 
signal s143	: std_logic_vector(31 downto 0); 
signal s144	: std_logic_vector(31 downto 0); 
signal s145	: std_logic_vector(31 downto 0); 
signal s147	: std_logic_vector(31 downto 0); 
signal s148	: std_logic_vector(31 downto 0); 
signal s373	: std_logic_vector(31 downto 0); 
signal s150	: std_logic_vector(31 downto 0); 
signal s151	: std_logic_vector(31 downto 0); 
signal s152	: std_logic_vector(31 downto 0); 
signal s154	: std_logic_vector(31 downto 0); 
signal s155	: std_logic_vector(31 downto 0); 
signal s374	: std_logic_vector(31 downto 0); 
signal s157	: std_logic_vector(31 downto 0); 
signal s158	: std_logic_vector(31 downto 0); 
signal s159	: std_logic_vector(31 downto 0); 
signal s161	: std_logic_vector(31 downto 0); 
signal s162	: std_logic_vector(31 downto 0); 
signal s375	: std_logic_vector(31 downto 0); 
signal s164	: std_logic_vector(31 downto 0); 
signal s165	: std_logic_vector(31 downto 0); 
signal s166	: std_logic_vector(31 downto 0); 
signal s168	: std_logic_vector(31 downto 0); 
signal s169	: std_logic_vector(31 downto 0); 
signal s376	: std_logic_vector(31 downto 0); 
signal s171	: std_logic_vector(31 downto 0); 
signal s172	: std_logic_vector(31 downto 0); 
signal s173	: std_logic_vector(31 downto 0); 
signal s175	: std_logic_vector(31 downto 0); 
signal s176	: std_logic_vector(31 downto 0); 
signal s377	: std_logic_vector(31 downto 0); 
signal s178	: std_logic_vector(31 downto 0); 
signal s179	: std_logic_vector(31 downto 0); 
signal s180	: std_logic_vector(31 downto 0); 
signal s182	: std_logic_vector(31 downto 0); 
signal s183	: std_logic_vector(31 downto 0); 
signal s378	: std_logic_vector(31 downto 0); 
signal s185	: std_logic_vector(31 downto 0); 
signal s186	: std_logic_vector(31 downto 0); 
signal s187	: std_logic_vector(31 downto 0); 
signal s189	: std_logic_vector(31 downto 0); 
signal s190	: std_logic_vector(31 downto 0); 
signal s379	: std_logic_vector(31 downto 0); 
signal s192	: std_logic_vector(31 downto 0); 
signal s193	: std_logic_vector(31 downto 0); 
signal s194	: std_logic_vector(31 downto 0); 
signal s196	: std_logic_vector(31 downto 0); 
signal s197	: std_logic_vector(31 downto 0); 
signal s380	: std_logic_vector(31 downto 0); 
signal s199	: std_logic_vector(31 downto 0); 
signal s200	: std_logic_vector(31 downto 0); 
signal s201	: std_logic_vector(31 downto 0); 
signal s203	: std_logic_vector(31 downto 0); 
signal s204	: std_logic_vector(31 downto 0); 
signal s381	: std_logic_vector(31 downto 0); 
signal s206	: std_logic_vector(31 downto 0); 
signal s207	: std_logic_vector(31 downto 0); 
signal s208	: std_logic_vector(31 downto 0); 
signal s210	: std_logic_vector(31 downto 0); 
signal s211	: std_logic_vector(31 downto 0); 
signal s382	: std_logic_vector(31 downto 0); 
signal s213	: std_logic_vector(31 downto 0); 
signal s214	: std_logic_vector(31 downto 0); 
signal s215	: std_logic_vector(31 downto 0); 
signal s217	: std_logic_vector(31 downto 0); 
signal s218	: std_logic_vector(31 downto 0); 
signal s383	: std_logic_vector(31 downto 0); 
signal s220	: std_logic_vector(31 downto 0); 
signal s221	: std_logic_vector(31 downto 0); 
signal s223	: std_logic_vector(31 downto 0); 
signal s225	: std_logic_vector(31 downto 0); 
signal s227	: std_logic_vector(31 downto 0); 
signal s229	: std_logic_vector(31 downto 0); 
signal s231	: std_logic_vector(31 downto 0); 
signal s233	: std_logic_vector(31 downto 0); 
signal s235	: std_logic_vector(31 downto 0); 
signal s237	: std_logic_vector(31 downto 0); 
signal s239	: std_logic_vector(31 downto 0); 
signal s241	: std_logic_vector(31 downto 0); 
signal s243	: std_logic_vector(31 downto 0); 
signal s245	: std_logic_vector(31 downto 0); 
signal s247	: std_logic_vector(31 downto 0); 
signal s249	: std_logic_vector(31 downto 0); 
signal s251	: std_logic_vector(31 downto 0); 
signal s253	: std_logic_vector(31 downto 0); 
signal s255	: std_logic_vector(31 downto 0); 
signal s257	: std_logic_vector(31 downto 0); 
signal s259	: std_logic_vector(31 downto 0); 
signal s261	: std_logic_vector(31 downto 0); 
signal s263	: std_logic_vector(31 downto 0); 
signal s265	: std_logic_vector(31 downto 0); 
signal s267	: std_logic_vector(31 downto 0); 
signal s269	: std_logic_vector(31 downto 0); 
signal s271	: std_logic_vector(31 downto 0); 
signal s273	: std_logic_vector(31 downto 0); 
signal s275	: std_logic_vector(31 downto 0); 
signal s277	: std_logic_vector(31 downto 0); 
signal s279	: std_logic_vector(31 downto 0); 
signal s281	: std_logic_vector(31 downto 0); 
signal s283	: std_logic_vector(31 downto 0); 
signal s285	: std_logic_vector(31 downto 0); 
signal s287	: std_logic; 
signal s350	: std_logic_vector(31 downto 0); 
signal s351	: std_logic_vector(31 downto 0); 
signal s384	: std_logic_vector(31 downto 0); 
signal s385	: std_logic_vector(31 downto 0); 
signal s386	: std_logic_vector(31 downto 0); 
signal s387	: std_logic_vector(31 downto 0); 
signal s388	: std_logic_vector(31 downto 0); 
signal s389	: std_logic_vector(31 downto 0); 
signal s390	: std_logic_vector(31 downto 0); 
signal s391	: std_logic_vector(31 downto 0); 
signal s392	: std_logic_vector(31 downto 0); 
signal s393	: std_logic_vector(31 downto 0); 
signal s394	: std_logic_vector(31 downto 0); 
signal s395	: std_logic_vector(31 downto 0); 
signal s396	: std_logic_vector(31 downto 0); 
signal s397	: std_logic_vector(31 downto 0); 
signal s398	: std_logic_vector(31 downto 0); 
signal s399	: std_logic_vector(31 downto 0); 
signal s400	: std_logic_vector(31 downto 0); 
signal s401	: std_logic_vector(31 downto 0); 
signal s402	: std_logic_vector(31 downto 0); 
signal s403	: std_logic_vector(31 downto 0); 
signal s404	: std_logic_vector(31 downto 0); 
signal s405	: std_logic_vector(31 downto 0); 
signal s406	: std_logic_vector(31 downto 0); 
signal s407	: std_logic_vector(31 downto 0); 
signal s408	: std_logic_vector(31 downto 0); 
signal s409	: std_logic_vector(31 downto 0); 
signal s410	: std_logic_vector(31 downto 0); 
signal s411	: std_logic_vector(31 downto 0); 
signal s412	: std_logic_vector(31 downto 0); 
signal s413	: std_logic_vector(31 downto 0); 
signal s414	: std_logic_vector(31 downto 0); 
signal s480	: std_logic_vector(0 downto 0); 
signal s447	: std_logic; 
signal s448	: std_logic; 
signal s449	: std_logic_vector(0 downto 0); 

begin 

	\i\: counter
	generic map ( 
		bits => 32,
		condition => 1,
		down => 0,
		increment => 32,
		steps => 1
	)
	port map ( 
		clk => \clk\,
		clk_en => s447,
		done => s448,
		input => s351,
		output => s216,
		reset => \reset\,
		step => s287,
		termination => s350
	);

	\x\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s216,
		O0 => s223,
		reset => \reset\,
		we => s287
	);

	\sum\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s352,
		I1 => s1,
		O0 => s352,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_mult_op_s_b\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s3,
		I1 => s4,
		O0 => s1
	);

	\a\: block_ram_a
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s223(10 downto 0),
		clk => \clk\,
		data_out => s3
	);

	\b\: block_ram_b
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s223(10 downto 0),
		clk => \clk\,
		data_out => s4
	);

	\x_13\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s5,
		O0 => s225,
		reset => \reset\,
		we => s287
	);

	\i_15_add_op_s_c15\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s7,
		O0 => s5
	);

	\sum_17\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s353,
		I1 => s8,
		O0 => s353,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_19_mult_op_s_b_20\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s10,
		I1 => s11,
		O0 => s8
	);

	\a_19\: block_ram_a_19
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s225(10 downto 0),
		clk => \clk\,
		data_out => s10
	);

	\b_20\: block_ram_b_20
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s225(10 downto 0),
		clk => \clk\,
		data_out => s11
	);

	\x_21\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s12,
		O0 => s227,
		reset => \reset\,
		we => s287
	);

	\i_23_add_op_s_c23\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s14,
		O0 => s12
	);

	\sum_25\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s354,
		I1 => s15,
		O0 => s354,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_27_mult_op_s_b_28\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s17,
		I1 => s18,
		O0 => s15
	);

	\a_27\: block_ram_a_27
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s227(10 downto 0),
		clk => \clk\,
		data_out => s17
	);

	\b_28\: block_ram_b_28
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s227(10 downto 0),
		clk => \clk\,
		data_out => s18
	);

	\x_29\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s19,
		O0 => s229,
		reset => \reset\,
		we => s287
	);

	\i_31_add_op_s_c31\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s21,
		O0 => s19
	);

	\sum_33\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s355,
		I1 => s22,
		O0 => s355,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_35_mult_op_s_b_36\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s24,
		I1 => s25,
		O0 => s22
	);

	\a_35\: block_ram_a_35
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s229(10 downto 0),
		clk => \clk\,
		data_out => s24
	);

	\b_36\: block_ram_b_36
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s229(10 downto 0),
		clk => \clk\,
		data_out => s25
	);

	\x_37\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s26,
		O0 => s231,
		reset => \reset\,
		we => s287
	);

	\i_39_add_op_s_c39\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s28,
		O0 => s26
	);

	\sum_41\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s356,
		I1 => s29,
		O0 => s356,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_43_mult_op_s_b_44\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s31,
		I1 => s32,
		O0 => s29
	);

	\a_43\: block_ram_a_43
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s231(10 downto 0),
		clk => \clk\,
		data_out => s31
	);

	\b_44\: block_ram_b_44
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s231(10 downto 0),
		clk => \clk\,
		data_out => s32
	);

	\x_45\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s33,
		O0 => s233,
		reset => \reset\,
		we => s287
	);

	\i_47_add_op_s_c47\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s35,
		O0 => s33
	);

	\sum_49\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s357,
		I1 => s36,
		O0 => s357,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_51_mult_op_s_b_52\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s38,
		I1 => s39,
		O0 => s36
	);

	\a_51\: block_ram_a_51
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s233(10 downto 0),
		clk => \clk\,
		data_out => s38
	);

	\b_52\: block_ram_b_52
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s233(10 downto 0),
		clk => \clk\,
		data_out => s39
	);

	\x_53\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s40,
		O0 => s235,
		reset => \reset\,
		we => s287
	);

	\i_55_add_op_s_c55\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s42,
		O0 => s40
	);

	\sum_57\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s358,
		I1 => s43,
		O0 => s358,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_59_mult_op_s_b_60\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s45,
		I1 => s46,
		O0 => s43
	);

	\a_59\: block_ram_a_59
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s235(10 downto 0),
		clk => \clk\,
		data_out => s45
	);

	\b_60\: block_ram_b_60
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s235(10 downto 0),
		clk => \clk\,
		data_out => s46
	);

	\x_61\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s47,
		O0 => s237,
		reset => \reset\,
		we => s287
	);

	\i_63_add_op_s_c63\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s49,
		O0 => s47
	);

	\sum_65\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s359,
		I1 => s50,
		O0 => s359,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_67_mult_op_s_b_68\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s52,
		I1 => s53,
		O0 => s50
	);

	\a_67\: block_ram_a_67
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s237(10 downto 0),
		clk => \clk\,
		data_out => s52
	);

	\b_68\: block_ram_b_68
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s237(10 downto 0),
		clk => \clk\,
		data_out => s53
	);

	\x_69\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s54,
		O0 => s239,
		reset => \reset\,
		we => s287
	);

	\i_71_add_op_s_c71\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s56,
		O0 => s54
	);

	\sum_73\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s360,
		I1 => s57,
		O0 => s360,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_75_mult_op_s_b_76\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s59,
		I1 => s60,
		O0 => s57
	);

	\a_75\: block_ram_a_75
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s239(10 downto 0),
		clk => \clk\,
		data_out => s59
	);

	\b_76\: block_ram_b_76
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s239(10 downto 0),
		clk => \clk\,
		data_out => s60
	);

	\x_77\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s61,
		O0 => s241,
		reset => \reset\,
		we => s287
	);

	\i_79_add_op_s_c79\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s63,
		O0 => s61
	);

	\sum_81\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s361,
		I1 => s64,
		O0 => s361,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_83_mult_op_s_b_84\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s66,
		I1 => s67,
		O0 => s64
	);

	\a_83\: block_ram_a_83
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s241(10 downto 0),
		clk => \clk\,
		data_out => s66
	);

	\b_84\: block_ram_b_84
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s241(10 downto 0),
		clk => \clk\,
		data_out => s67
	);

	\x_85\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s68,
		O0 => s243,
		reset => \reset\,
		we => s287
	);

	\i_87_add_op_s_c87\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s70,
		O0 => s68
	);

	\sum_89\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s362,
		I1 => s71,
		O0 => s362,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_91_mult_op_s_b_92\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s73,
		I1 => s74,
		O0 => s71
	);

	\a_91\: block_ram_a_91
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s243(10 downto 0),
		clk => \clk\,
		data_out => s73
	);

	\b_92\: block_ram_b_92
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s243(10 downto 0),
		clk => \clk\,
		data_out => s74
	);

	\x_93\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s75,
		O0 => s245,
		reset => \reset\,
		we => s287
	);

	\i_95_add_op_s_c95\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s77,
		O0 => s75
	);

	\sum_97\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s363,
		I1 => s78,
		O0 => s363,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_99_mult_op_s_b_100\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s80,
		I1 => s81,
		O0 => s78
	);

	\a_99\: block_ram_a_99
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s245(10 downto 0),
		clk => \clk\,
		data_out => s80
	);

	\b_100\: block_ram_b_100
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s245(10 downto 0),
		clk => \clk\,
		data_out => s81
	);

	\x_101\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s82,
		O0 => s247,
		reset => \reset\,
		we => s287
	);

	\i_103_add_op_s_c103\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s84,
		O0 => s82
	);

	\sum_105\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s364,
		I1 => s85,
		O0 => s364,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_107_mult_op_s_b_108\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s87,
		I1 => s88,
		O0 => s85
	);

	\a_107\: block_ram_a_107
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s247(10 downto 0),
		clk => \clk\,
		data_out => s87
	);

	\b_108\: block_ram_b_108
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s247(10 downto 0),
		clk => \clk\,
		data_out => s88
	);

	\x_109\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s89,
		O0 => s249,
		reset => \reset\,
		we => s287
	);

	\i_111_add_op_s_c111\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s91,
		O0 => s89
	);

	\sum_113\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s365,
		I1 => s92,
		O0 => s365,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_115_mult_op_s_b_116\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s94,
		I1 => s95,
		O0 => s92
	);

	\a_115\: block_ram_a_115
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s249(10 downto 0),
		clk => \clk\,
		data_out => s94
	);

	\b_116\: block_ram_b_116
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s249(10 downto 0),
		clk => \clk\,
		data_out => s95
	);

	\x_117\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s96,
		O0 => s251,
		reset => \reset\,
		we => s287
	);

	\i_119_add_op_s_c119\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s98,
		O0 => s96
	);

	\sum_121\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s366,
		I1 => s99,
		O0 => s366,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_123_mult_op_s_b_124\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s101,
		I1 => s102,
		O0 => s99
	);

	\a_123\: block_ram_a_123
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s251(10 downto 0),
		clk => \clk\,
		data_out => s101
	);

	\b_124\: block_ram_b_124
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s251(10 downto 0),
		clk => \clk\,
		data_out => s102
	);

	\x_125\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s103,
		O0 => s253,
		reset => \reset\,
		we => s287
	);

	\i_127_add_op_s_c127\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s105,
		O0 => s103
	);

	\sum_129\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s367,
		I1 => s106,
		O0 => s367,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_131_mult_op_s_b_132\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s108,
		I1 => s109,
		O0 => s106
	);

	\a_131\: block_ram_a_131
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s253(10 downto 0),
		clk => \clk\,
		data_out => s108
	);

	\b_132\: block_ram_b_132
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s253(10 downto 0),
		clk => \clk\,
		data_out => s109
	);

	\x_133\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s110,
		O0 => s255,
		reset => \reset\,
		we => s287
	);

	\i_135_add_op_s_c135\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s112,
		O0 => s110
	);

	\sum_137\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s368,
		I1 => s113,
		O0 => s368,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_139_mult_op_s_b_140\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s115,
		I1 => s116,
		O0 => s113
	);

	\a_139\: block_ram_a_139
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s255(10 downto 0),
		clk => \clk\,
		data_out => s115
	);

	\b_140\: block_ram_b_140
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s255(10 downto 0),
		clk => \clk\,
		data_out => s116
	);

	\x_141\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s117,
		O0 => s257,
		reset => \reset\,
		we => s287
	);

	\i_143_add_op_s_c143\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s119,
		O0 => s117
	);

	\sum_145\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s369,
		I1 => s120,
		O0 => s369,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_147_mult_op_s_b_148\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s122,
		I1 => s123,
		O0 => s120
	);

	\a_147\: block_ram_a_147
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s257(10 downto 0),
		clk => \clk\,
		data_out => s122
	);

	\b_148\: block_ram_b_148
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s257(10 downto 0),
		clk => \clk\,
		data_out => s123
	);

	\x_149\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s124,
		O0 => s259,
		reset => \reset\,
		we => s287
	);

	\i_151_add_op_s_c151\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s126,
		O0 => s124
	);

	\sum_153\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s370,
		I1 => s127,
		O0 => s370,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_155_mult_op_s_b_156\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s129,
		I1 => s130,
		O0 => s127
	);

	\a_155\: block_ram_a_155
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s259(10 downto 0),
		clk => \clk\,
		data_out => s129
	);

	\b_156\: block_ram_b_156
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s259(10 downto 0),
		clk => \clk\,
		data_out => s130
	);

	\x_157\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s131,
		O0 => s261,
		reset => \reset\,
		we => s287
	);

	\i_159_add_op_s_c159\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s133,
		O0 => s131
	);

	\sum_161\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s371,
		I1 => s134,
		O0 => s371,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_163_mult_op_s_b_164\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s136,
		I1 => s137,
		O0 => s134
	);

	\a_163\: block_ram_a_163
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s261(10 downto 0),
		clk => \clk\,
		data_out => s136
	);

	\b_164\: block_ram_b_164
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s261(10 downto 0),
		clk => \clk\,
		data_out => s137
	);

	\x_165\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s138,
		O0 => s263,
		reset => \reset\,
		we => s287
	);

	\i_167_add_op_s_c167\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s140,
		O0 => s138
	);

	\sum_169\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s372,
		I1 => s141,
		O0 => s372,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_171_mult_op_s_b_172\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s143,
		I1 => s144,
		O0 => s141
	);

	\a_171\: block_ram_a_171
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s263(10 downto 0),
		clk => \clk\,
		data_out => s143
	);

	\b_172\: block_ram_b_172
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s263(10 downto 0),
		clk => \clk\,
		data_out => s144
	);

	\x_173\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s145,
		O0 => s265,
		reset => \reset\,
		we => s287
	);

	\i_175_add_op_s_c175\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s147,
		O0 => s145
	);

	\sum_177\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s373,
		I1 => s148,
		O0 => s373,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_179_mult_op_s_b_180\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s150,
		I1 => s151,
		O0 => s148
	);

	\a_179\: block_ram_a_179
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s265(10 downto 0),
		clk => \clk\,
		data_out => s150
	);

	\b_180\: block_ram_b_180
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s265(10 downto 0),
		clk => \clk\,
		data_out => s151
	);

	\x_181\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s152,
		O0 => s267,
		reset => \reset\,
		we => s287
	);

	\i_183_add_op_s_c183\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s154,
		O0 => s152
	);

	\sum_185\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s374,
		I1 => s155,
		O0 => s374,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_187_mult_op_s_b_188\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s157,
		I1 => s158,
		O0 => s155
	);

	\a_187\: block_ram_a_187
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s267(10 downto 0),
		clk => \clk\,
		data_out => s157
	);

	\b_188\: block_ram_b_188
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s267(10 downto 0),
		clk => \clk\,
		data_out => s158
	);

	\x_189\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s159,
		O0 => s269,
		reset => \reset\,
		we => s287
	);

	\i_191_add_op_s_c191\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s161,
		O0 => s159
	);

	\sum_193\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s375,
		I1 => s162,
		O0 => s375,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_195_mult_op_s_b_196\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s164,
		I1 => s165,
		O0 => s162
	);

	\a_195\: block_ram_a_195
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s269(10 downto 0),
		clk => \clk\,
		data_out => s164
	);

	\b_196\: block_ram_b_196
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s269(10 downto 0),
		clk => \clk\,
		data_out => s165
	);

	\x_197\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s166,
		O0 => s271,
		reset => \reset\,
		we => s287
	);

	\i_199_add_op_s_c199\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s168,
		O0 => s166
	);

	\sum_201\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s376,
		I1 => s169,
		O0 => s376,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_203_mult_op_s_b_204\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s171,
		I1 => s172,
		O0 => s169
	);

	\a_203\: block_ram_a_203
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s271(10 downto 0),
		clk => \clk\,
		data_out => s171
	);

	\b_204\: block_ram_b_204
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s271(10 downto 0),
		clk => \clk\,
		data_out => s172
	);

	\x_205\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s173,
		O0 => s273,
		reset => \reset\,
		we => s287
	);

	\i_207_add_op_s_c207\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s175,
		O0 => s173
	);

	\sum_209\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s377,
		I1 => s176,
		O0 => s377,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_211_mult_op_s_b_212\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s178,
		I1 => s179,
		O0 => s176
	);

	\a_211\: block_ram_a_211
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s273(10 downto 0),
		clk => \clk\,
		data_out => s178
	);

	\b_212\: block_ram_b_212
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s273(10 downto 0),
		clk => \clk\,
		data_out => s179
	);

	\x_213\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s180,
		O0 => s275,
		reset => \reset\,
		we => s287
	);

	\i_215_add_op_s_c215\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s182,
		O0 => s180
	);

	\sum_217\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s378,
		I1 => s183,
		O0 => s378,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_219_mult_op_s_b_220\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s185,
		I1 => s186,
		O0 => s183
	);

	\a_219\: block_ram_a_219
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s275(10 downto 0),
		clk => \clk\,
		data_out => s185
	);

	\b_220\: block_ram_b_220
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s275(10 downto 0),
		clk => \clk\,
		data_out => s186
	);

	\x_221\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s187,
		O0 => s277,
		reset => \reset\,
		we => s287
	);

	\i_223_add_op_s_c223\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s189,
		O0 => s187
	);

	\sum_225\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s379,
		I1 => s190,
		O0 => s379,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_227_mult_op_s_b_228\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s192,
		I1 => s193,
		O0 => s190
	);

	\a_227\: block_ram_a_227
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s277(10 downto 0),
		clk => \clk\,
		data_out => s192
	);

	\b_228\: block_ram_b_228
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s277(10 downto 0),
		clk => \clk\,
		data_out => s193
	);

	\x_229\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s194,
		O0 => s279,
		reset => \reset\,
		we => s287
	);

	\i_231_add_op_s_c231\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s196,
		O0 => s194
	);

	\sum_233\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s380,
		I1 => s197,
		O0 => s380,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_235_mult_op_s_b_236\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s199,
		I1 => s200,
		O0 => s197
	);

	\a_235\: block_ram_a_235
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s279(10 downto 0),
		clk => \clk\,
		data_out => s199
	);

	\b_236\: block_ram_b_236
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s279(10 downto 0),
		clk => \clk\,
		data_out => s200
	);

	\x_237\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s201,
		O0 => s281,
		reset => \reset\,
		we => s287
	);

	\i_239_add_op_s_c239\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s203,
		O0 => s201
	);

	\sum_241\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s381,
		I1 => s204,
		O0 => s381,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_243_mult_op_s_b_244\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s206,
		I1 => s207,
		O0 => s204
	);

	\a_243\: block_ram_a_243
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s281(10 downto 0),
		clk => \clk\,
		data_out => s206
	);

	\b_244\: block_ram_b_244
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s281(10 downto 0),
		clk => \clk\,
		data_out => s207
	);

	\x_245\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s208,
		O0 => s283,
		reset => \reset\,
		we => s287
	);

	\i_247_add_op_s_c247\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s210,
		O0 => s208
	);

	\sum_249\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s382,
		I1 => s211,
		O0 => s382,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_251_mult_op_s_b_252\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s213,
		I1 => s214,
		O0 => s211
	);

	\a_251\: block_ram_a_251
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s283(10 downto 0),
		clk => \clk\,
		data_out => s213
	);

	\b_252\: block_ram_b_252
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s283(10 downto 0),
		clk => \clk\,
		data_out => s214
	);

	\x_253\: reg_op
	generic map ( 
		initial => 0,
		w_in => 32
	)
	port map ( 
		clk => \clk\,
		I0 => s215,
		O0 => s285,
		reset => \reset\,
		we => s287
	);

	\i_255_add_op_s_c255\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s216,
		I1 => s217,
		O0 => s215
	);

	\sum_257\: add_reg_op_s
	generic map ( 
		initial => 0,
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s383,
		I1 => s218,
		O0 => s383,
		clk => \clk\,
		reset => \reset\,
		we => s480(0)
	);

	\a_259_mult_op_s_b_260\: mult_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s220,
		I1 => s221,
		O0 => s218
	);

	\a_259\: block_ram_a_259
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s285(10 downto 0),
		clk => \clk\,
		data_out => s220
	);

	\b_260\: block_ram_b_260
	generic map ( 
		address_width => 11,
		data_width => 32
	)
	port map ( 
		address(10 downto 0) => s285(10 downto 0),
		clk => \clk\,
		data_out => s221
	);

	\sum_add_op_s_sum_17\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s352,
		I1 => s353,
		O0 => s384
	);

	\sum_25_add_op_s_sum_33\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s354,
		I1 => s355,
		O0 => s385
	);

	\sum_41_add_op_s_sum_49\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s356,
		I1 => s357,
		O0 => s386
	);

	\sum_57_add_op_s_sum_65\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s358,
		I1 => s359,
		O0 => s387
	);

	\sum_73_add_op_s_sum_81\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s360,
		I1 => s361,
		O0 => s388
	);

	\sum_89_add_op_s_sum_97\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s362,
		I1 => s363,
		O0 => s389
	);

	\sum_105_add_op_s_sum_113\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s364,
		I1 => s365,
		O0 => s390
	);

	\sum_121_add_op_s_sum_129\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s366,
		I1 => s367,
		O0 => s391
	);

	\sum_137_add_op_s_sum_145\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s368,
		I1 => s369,
		O0 => s392
	);

	\sum_153_add_op_s_sum_161\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s370,
		I1 => s371,
		O0 => s393
	);

	\sum_169_add_op_s_sum_177\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s372,
		I1 => s373,
		O0 => s394
	);

	\sum_185_add_op_s_sum_193\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s374,
		I1 => s375,
		O0 => s395
	);

	\sum_201_add_op_s_sum_209\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s376,
		I1 => s377,
		O0 => s396
	);

	\sum_217_add_op_s_sum_225\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s378,
		I1 => s379,
		O0 => s397
	);

	\sum_233_add_op_s_sum_241\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s380,
		I1 => s381,
		O0 => s398
	);

	\sum_249_add_op_s_sum_257\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s382,
		I1 => s383,
		O0 => s399
	);

	\sum_add_op_s_sum_17_add_op_s_sum_25_add_op_s_sum_33\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s384,
		I1 => s385,
		O0 => s400
	);

	\sum_41_add_op_s_sum_49_add_op_s_sum_57_add_op_s_sum_65\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s386,
		I1 => s387,
		O0 => s401
	);

	\sum_73_add_op_s_sum_81_add_op_s_sum_89_add_op_s_sum_97\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s388,
		I1 => s389,
		O0 => s402
	);

	\sum_105_add_op_s_sum_113_add_op_s_sum_121_add_op_s_sum_129\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s390,
		I1 => s391,
		O0 => s403
	);

	\sum_137_add_op_s_sum_145_add_op_s_sum_153_add_op_s_sum_161\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s392,
		I1 => s393,
		O0 => s404
	);

	\sum_169_add_op_s_sum_177_add_op_s_sum_185_add_op_s_sum_193\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s394,
		I1 => s395,
		O0 => s405
	);

	\sum_201_add_op_s_sum_209_add_op_s_sum_217_add_op_s_sum_225\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s396,
		I1 => s397,
		O0 => s406
	);

	\sum_233_add_op_s_sum_241_add_op_s_sum_249_add_op_s_sum_257\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s398,
		I1 => s399,
		O0 => s407
	);

	\sum_add_op_s_sum_17_add_op_s_sum_25_add_op_s_sum_33_add_op_s_sum_41_add_op_s_sum_49_add_op_s_sum_57_add_op_s_sum_65\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s400,
		I1 => s401,
		O0 => s408
	);

	\sum_73_add_op_s_sum_81_add_op_s_sum_89_add_op_s_sum_97_add_op_s_sum_105_add_op_s_sum_113_add_op_s_sum_121_add_op_s_sum_129\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s402,
		I1 => s403,
		O0 => s409
	);

	\sum_137_add_op_s_sum_145_add_op_s_sum_153_add_op_s_sum_161_add_op_s_sum_169_add_op_s_sum_177_add_op_s_sum_185_add_op_s_sum_193\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s404,
		I1 => s405,
		O0 => s410
	);

	\sum_201_add_op_s_sum_209_add_op_s_sum_217_add_op_s_sum_225_add_op_s_sum_233_add_op_s_sum_241_add_op_s_sum_249_add_op_s_sum_257\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s406,
		I1 => s407,
		O0 => s411
	);

	\sum_add_op_s_sum_17_add_op_s_sum_25_add_op_s_sum_33_add_op_s_sum_41_add_op_s_sum_49_add_op_s_sum_57_add_op_s_sum_65_add_op_s_sum_73_add_op_s_sum_81_add_op_s_sum_89_add_op_s_sum_97_add_op_s_sum_105_add_op_s_sum_113_add_op_s_sum_121_add_op_s_sum_129\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s408,
		I1 => s409,
		O0 => s412
	);

	\sum_137_add_op_s_sum_145_add_op_s_sum_153_add_op_s_sum_161_add_op_s_sum_169_add_op_s_sum_177_add_op_s_sum_185_add_op_s_sum_193_add_op_s_sum_201_add_op_s_sum_209_add_op_s_sum_217_add_op_s_sum_225_add_op_s_sum_233_add_op_s_sum_241_add_op_s_sum_249_add_op_s_sum_257\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s410,
		I1 => s411,
		O0 => s413
	);

	\sum_add_op_s_sum_17_add_op_s_sum_25_add_op_s_sum_33_add_op_s_sum_41_add_op_s_sum_49_add_op_s_sum_57_add_op_s_sum_65_add_op_s_sum_73_add_op_s_sum_81_add_op_s_sum_89_add_op_s_sum_97_add_op_s_sum_105_add_op_s_sum_113_add_op_s_sum_121_add_op_s_sum_129_add_op_s_sum_137_add_op_s_sum_145_add_op_s_sum_153_add_op_s_sum_161_add_op_s_sum_169_add_op_s_sum_177_add_op_s_sum_185_add_op_s_sum_193_add_op_s_sum_201_add_op_s_sum_209_add_op_s_sum_217_add_op_s_sum_225_add_op_s_sum_233_add_op_s_sum_241_add_op_s_sum_249_add_op_s_sum_257\: add_op_s
	generic map ( 
		w_in1 => 32,
		w_in2 => 32,
		w_out => 32
	)
	port map ( 
		I0 => s412,
		I1 => s413,
		O0 => s414
	);

	\c420\: delay_op
	generic map ( 
		bits => 1,
		delay => 3
	)
	port map ( 
		a(0) => s287,
		a_delayed => s480,
		clk => \clk\,
		reset => \reset\
	);

	\c452\: delay_op
	generic map ( 
		bits => 1,
		delay => 7
	)
	port map ( 
		a(0) => s448,
		a_delayed => s449,
		clk => \clk\,
		reset => \reset\
	);

s7 <= conv_std_logic_vector(1, 32); 
s14 <= conv_std_logic_vector(2, 32); 
s21 <= conv_std_logic_vector(3, 32); 
s28 <= conv_std_logic_vector(4, 32); 
s35 <= conv_std_logic_vector(5, 32); 
s42 <= conv_std_logic_vector(6, 32); 
s49 <= conv_std_logic_vector(7, 32); 
s56 <= conv_std_logic_vector(8, 32); 
s63 <= conv_std_logic_vector(9, 32); 
s70 <= conv_std_logic_vector(10, 32); 
s77 <= conv_std_logic_vector(11, 32); 
s84 <= conv_std_logic_vector(12, 32); 
s91 <= conv_std_logic_vector(13, 32); 
s98 <= conv_std_logic_vector(14, 32); 
s105 <= conv_std_logic_vector(15, 32); 
s112 <= conv_std_logic_vector(16, 32); 
s119 <= conv_std_logic_vector(17, 32); 
s126 <= conv_std_logic_vector(18, 32); 
s133 <= conv_std_logic_vector(19, 32); 
s140 <= conv_std_logic_vector(20, 32); 
s147 <= conv_std_logic_vector(21, 32); 
s154 <= conv_std_logic_vector(22, 32); 
s161 <= conv_std_logic_vector(23, 32); 
s168 <= conv_std_logic_vector(24, 32); 
s175 <= conv_std_logic_vector(25, 32); 
s182 <= conv_std_logic_vector(26, 32); 
s189 <= conv_std_logic_vector(27, 32); 
s196 <= conv_std_logic_vector(28, 32); 
s203 <= conv_std_logic_vector(29, 32); 
s210 <= conv_std_logic_vector(30, 32); 
s217 <= conv_std_logic_vector(31, 32); 
s447 <= \init\; 
\done\ <= s449(0); 
s350 <= conv_std_logic_vector(2047, 32); 
s351 <= conv_std_logic_vector(0, 32); 
\result\ <= s414; 
end behavior; 