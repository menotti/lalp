library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 
entity sobel_multport_f2 is 
	port (
		\init\	: in	std_logic;
		\done\	: out	std_logic;
		\out_257\	: out	std_logic_vector(31 downto 0);
		\out_258\	: out	std_logic_vector(31 downto 0);
		\clk\	: in	std_logic;
		\reset\	: in	std_logic;
		\clear\	: in	std_logic
	);
end sobel_multport_f2; 

architecture behavior of sobel_multport_f2 is 

component add_op_s 
generic ( 
        w_in1	: integer := 8; 
        w_in2	: integer := 8; 
        w_out	: integer := 16 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component block_ram_mult_in 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        address_0           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_0           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_0          :out    std_logic_vector (data_width-1 downto 0); 
        we_0                :in     std_logic := '0'; 
        oe_0                :in     std_logic := '1'; 
        address_1           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_1           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_1          :out    std_logic_vector (data_width-1 downto 0); 
        we_1                :in     std_logic := '0'; 
        oe_1                :in     std_logic := '1'; 
        address_2           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_2           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_2          :out    std_logic_vector (data_width-1 downto 0); 
        we_2                :in     std_logic := '0'; 
        oe_2                :in     std_logic := '1'; 
        address_3           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_3           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_3          :out    std_logic_vector (data_width-1 downto 0); 
        we_3                :in     std_logic := '0'; 
        oe_3                :in     std_logic := '1'; 
        address_4           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_4           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_4          :out    std_logic_vector (data_width-1 downto 0); 
        we_4                :in     std_logic := '0'; 
        oe_4                :in     std_logic := '1'; 
        address_5           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_5           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_5          :out    std_logic_vector (data_width-1 downto 0); 
        we_5                :in     std_logic := '0'; 
        oe_5                :in     std_logic := '1'; 
        address_6           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_6           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_6          :out    std_logic_vector (data_width-1 downto 0); 
        we_6                :in     std_logic := '0'; 
        oe_6                :in     std_logic := '1'; 
        address_7           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_7           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_7          :out    std_logic_vector (data_width-1 downto 0); 
        we_7                :in     std_logic := '0'; 
        oe_7                :in     std_logic := '1'; 
        address_8           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_8           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_8          :out    std_logic_vector (data_width-1 downto 0); 
        we_8                :in     std_logic := '0'; 
        oe_8                :in     std_logic := '1'; 
        address_9           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_9           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_9          :out    std_logic_vector (data_width-1 downto 0); 
        we_9                :in     std_logic := '0'; 
        oe_9                :in     std_logic := '1'; 
        address_10           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_10           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_10          :out    std_logic_vector (data_width-1 downto 0); 
        we_10                :in     std_logic := '0'; 
        oe_10                :in     std_logic := '1'; 
        address_11           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_11           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_11          :out    std_logic_vector (data_width-1 downto 0); 
        we_11                :in     std_logic := '0'; 
        oe_11                :in     std_logic := '1'; 
        address_12           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_12           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_12          :out    std_logic_vector (data_width-1 downto 0); 
        we_12                :in     std_logic := '0'; 
        oe_12                :in     std_logic := '1'; 
        address_13           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_13           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_13          :out    std_logic_vector (data_width-1 downto 0); 
        we_13                :in     std_logic := '0'; 
        oe_13                :in     std_logic := '1'; 
        address_14           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_14           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_14          :out    std_logic_vector (data_width-1 downto 0); 
        we_14                :in     std_logic := '0'; 
        oe_14                :in     std_logic := '1'; 
        address_15           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_15           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_15          :out    std_logic_vector (data_width-1 downto 0); 
        we_15                :in     std_logic := '0'; 
        oe_15                :in     std_logic := '1'; 
        clk                 :       in std_logic 
); 
end component; 

component block_ram_mult_out 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        address_0           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_0           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_0          :out    std_logic_vector (data_width-1 downto 0); 
        we_0                :in     std_logic := '0'; 
        oe_0                :in     std_logic := '1'; 
        address_1           :in     std_logic_vector (address_width-1 downto 0); 
        data_in_1           :in     std_logic_vector (data_width-1 downto 0) := (others => '0'); 
        data_out_1          :out    std_logic_vector (data_width-1 downto 0); 
        we_1                :in     std_logic := '0'; 
        oe_1                :in     std_logic := '1'; 
        clk                 :       in std_logic 
); 
end component; 

component counter 
generic (
        bits		: integer := 8;
        steps		: integer := 1;
        increment           : integer := 1;
        down                : integer := 0;
        condition           : integer := 0
);
port (
        input		: in	std_logic_vector(bits-1 downto 0);
        termination         : in	std_logic_vector(bits-1 downto 0);
        clk                 : in	std_logic;
        clk_en		: in	std_logic := '1';
        reset		: in	std_logic;
        load		: in	std_logic := '0';
        step		: out	std_logic;
        done		: out	std_logic;
        output		: out	std_logic_vector(bits-1 downto 0)
); 
end component; 

component delay_op 
generic ( 
        bits        : integer := 8; 
        delay       : integer := 1 
); 
port ( 
        a		: in	std_logic_vector(bits-1 downto 0); 
        clk		: in	std_logic; 
        reset	: in	std_logic; 
        a_delayed	: out	std_logic_vector(bits-1 downto 0) := (others=>'0') 
); 
end component; 

component if_gt_op_s 
generic ( 
        w_in1	: integer := 16; 
        w_in2	: integer := 16; 
        w_out	: integer := 1 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component if_lt_op_s 
generic ( 
        w_in1	: integer := 16; 
        w_in2	: integer := 16; 
        w_out	: integer := 1 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component neg_op_s 
generic ( 
        w_in        : integer := 16;
        w_out       : integer := 16 
); 
port ( 
        I0		: in	std_logic_vector(w_in-1 downto 0); 
        O0		: out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component reg_mux_op 
generic ( 
        w_in	: integer := 16; 
        initial	: integer := 0 
); 
port ( 
        clk         : in	std_logic; 
        reset       : in	std_logic; 
        we          : in	std_logic := '1'; 
        Sel1	: in	std_logic_vector(0 downto 0);
        I0          : in	std_logic_vector(w_in-1 downto 0); 
        I1          : in	std_logic_vector(w_in-1 downto 0); 
        O0          : out	std_logic_vector(w_in-1 downto 0) 
); 
end component; 

component reg_op 
generic ( 
        w_in	: integer := 16; 
        initial	: integer := 0 
); 
port ( 
        clk         : in	std_logic; 
        reset       : in	std_logic; 
        we          : in	std_logic := '1'; 
        I0          : in	std_logic_vector(w_in-1 downto 0); 
        O0          : out	std_logic_vector(w_in-1 downto 0) 
); 
end component; 

component sub_op_s 
generic ( 
        w_in1	: integer := 8; 
        w_in2	: integer := 8; 
        w_out	: integer := 16 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

signal s9	: std_logic_vector(31 downto 0); 
signal s11	: std_logic_vector(31 downto 0); 
signal s13	: std_logic_vector(31 downto 0); 
signal s24	: std_logic_vector(31 downto 0); 
signal s26	: std_logic_vector(31 downto 0); 
signal s28	: std_logic_vector(31 downto 0); 
signal s33	: std_logic_vector(31 downto 0); 
signal s36	: std_logic_vector(31 downto 0); 
signal s39	: std_logic_vector(31 downto 0); 
signal s42	: std_logic_vector(31 downto 0); 
signal s45	: std_logic_vector(31 downto 0); 
signal s48	: std_logic_vector(31 downto 0); 
signal s51	: std_logic_vector(31 downto 0); 
signal s52	: std_logic_vector(31 downto 0); 
signal s53	: std_logic_vector(31 downto 0); 
signal s54	: std_logic_vector(31 downto 0); 
signal s56	: std_logic_vector(31 downto 0); 
signal s57	: std_logic_vector(31 downto 0); 
signal s60	: std_logic_vector(31 downto 0); 
signal s61	: std_logic_vector(31 downto 0); 
signal s62	: std_logic_vector(31 downto 0); 
signal s65	: std_logic_vector(31 downto 0); 
signal s66	: std_logic_vector(31 downto 0); 
signal s70	: std_logic_vector(31 downto 0); 
signal s71	: std_logic_vector(31 downto 0); 
signal s72	: std_logic_vector(31 downto 0); 
signal s75	: std_logic_vector(31 downto 0); 
signal s76	: std_logic_vector(31 downto 0); 
signal s77	: std_logic_vector(31 downto 0); 
signal s78	: std_logic_vector(31 downto 0); 
signal s81	: std_logic_vector(31 downto 0); 
signal s84	: std_logic_vector(31 downto 0); 
signal s85	: std_logic_vector(31 downto 0); 
signal s92	: std_logic_vector(31 downto 0); 
signal s106	: std_logic_vector(31 downto 0); 
signal s108	: std_logic_vector(31 downto 0); 
signal s110	: std_logic_vector(31 downto 0); 
signal s112	: std_logic_vector(31 downto 0); 
signal s114	: std_logic_vector(31 downto 0); 
signal s116	: std_logic_vector(31 downto 0); 
signal s118	: std_logic_vector(31 downto 0); 
signal s120	: std_logic_vector(31 downto 0); 
signal s121	: std_logic_vector(31 downto 0); 
signal s122	: std_logic_vector(31 downto 0); 
signal s123	: std_logic_vector(31 downto 0); 
signal s125	: std_logic_vector(31 downto 0); 
signal s126	: std_logic_vector(31 downto 0); 
signal s129	: std_logic_vector(31 downto 0); 
signal s130	: std_logic_vector(31 downto 0); 
signal s131	: std_logic_vector(31 downto 0); 
signal s134	: std_logic_vector(31 downto 0); 
signal s135	: std_logic_vector(31 downto 0); 
signal s139	: std_logic_vector(31 downto 0); 
signal s140	: std_logic_vector(31 downto 0); 
signal s141	: std_logic_vector(31 downto 0); 
signal s144	: std_logic_vector(31 downto 0); 
signal s145	: std_logic_vector(31 downto 0); 
signal s146	: std_logic_vector(31 downto 0); 
signal s147	: std_logic_vector(31 downto 0); 
signal s150	: std_logic_vector(31 downto 0); 
signal s153	: std_logic_vector(31 downto 0); 
signal s154	: std_logic_vector(31 downto 0); 
signal s161	: std_logic_vector(31 downto 0); 
signal s166	: std_logic_vector(31 downto 0); 
signal s168	: std_logic_vector(0 downto 0); 
signal s169	: std_logic_vector(31 downto 0); 
signal s171	: std_logic_vector(0 downto 0); 
signal s172	: std_logic_vector(31 downto 0); 
signal s174	: std_logic_vector(0 downto 0); 
signal s175	: std_logic_vector(31 downto 0); 
signal s177	: std_logic_vector(0 downto 0); 
signal s178	: std_logic_vector(31 downto 0); 
signal s180	: std_logic_vector(0 downto 0); 
signal s181	: std_logic_vector(31 downto 0); 
signal s183	: std_logic_vector(0 downto 0); 
signal s185	: std_logic_vector(31 downto 0); 
signal s187	: std_logic_vector(31 downto 0); 
signal s189	: std_logic_vector(31 downto 0); 
signal s191	: std_logic_vector(31 downto 0); 
signal s193	: std_logic_vector(31 downto 0); 
signal s195	: std_logic_vector(31 downto 0); 
signal s197	: std_logic_vector(31 downto 0); 
signal s199	: std_logic_vector(31 downto 0); 
signal s201	: std_logic_vector(31 downto 0); 
signal s202	: std_logic_vector(31 downto 0); 
signal s204	: std_logic_vector(31 downto 0); 
signal s205	: std_logic_vector(31 downto 0); 
signal s206	: std_logic_vector(31 downto 0); 
signal s209	: std_logic_vector(31 downto 0); 
signal s211	: std_logic_vector(31 downto 0); 
signal s213	: std_logic_vector(31 downto 0); 
signal s215	: std_logic_vector(31 downto 0); 
signal s217	: std_logic_vector(31 downto 0); 
signal s219	: std_logic_vector(31 downto 0); 
signal s221	: std_logic_vector(31 downto 0); 
signal s223	: std_logic_vector(31 downto 0); 
signal s225	: std_logic_vector(31 downto 0); 
signal s226	: std_logic_vector(31 downto 0); 
signal s228	: std_logic_vector(31 downto 0); 
signal s229	: std_logic_vector(31 downto 0); 
signal s230	: std_logic_vector(31 downto 0); 
signal s232	: std_logic_vector(31 downto 0); 
signal s233	: std_logic_vector(31 downto 0); 
signal s238	: std_logic_vector(0 downto 0); 
signal s240	: std_logic_vector(0 downto 0); 
signal s242	: std_logic_vector(0 downto 0); 
signal s244	: std_logic_vector(0 downto 0); 
signal s246	: std_logic_vector(0 downto 0); 
signal s248	: std_logic_vector(0 downto 0); 
signal s250	: std_logic_vector(0 downto 0); 
signal s252	: std_logic_vector(0 downto 0); 
signal s254	: std_logic_vector(0 downto 0); 
signal s256	: std_logic_vector(0 downto 0); 
signal s258	: std_logic_vector(0 downto 0); 
signal s260	: std_logic_vector(0 downto 0); 
signal s262	: std_logic_vector(0 downto 0); 
signal s264	: std_logic_vector(0 downto 0); 
signal s266	: std_logic_vector(0 downto 0); 
signal s268	: std_logic_vector(0 downto 0); 
signal s270	: std_logic_vector(0 downto 0); 
signal s272	: std_logic_vector(0 downto 0); 
signal s274	: std_logic_vector(0 downto 0); 
signal s276	: std_logic_vector(0 downto 0); 
signal s278	: std_logic_vector(0 downto 0); 
signal s280	: std_logic_vector(0 downto 0); 
signal s282	: std_logic_vector(0 downto 0); 
signal s284	: std_logic_vector(0 downto 0); 
signal s286	: std_logic_vector(0 downto 0); 
signal s288	: std_logic_vector(0 downto 0); 
signal s290	: std_logic_vector(0 downto 0); 
signal s291	: std_logic; 
signal s292	: std_logic_vector(0 downto 0); 
signal s293	: std_logic; 
signal s294	: std_logic; 
signal s295	: std_logic_vector(0 downto 0); 
signal s299	: std_logic_vector(31 downto 0); 
signal s300	: std_logic_vector(31 downto 0); 
signal s301	: std_logic_vector(31 downto 0); 
signal s302	: std_logic_vector(31 downto 0); 
signal s303	: std_logic_vector(31 downto 0); 
signal s304	: std_logic_vector(31 downto 0); 
signal s305	: std_logic_vector(31 downto 0); 
signal s306	: std_logic_vector(31 downto 0); 
signal s307	: std_logic_vector(31 downto 0); 
signal s308	: std_logic_vector(31 downto 0); 
signal s309	: std_logic_vector(31 downto 0); 
signal s310	: std_logic_vector(31 downto 0); 
signal s311	: std_logic_vector(31 downto 0); 
signal s312	: std_logic_vector(31 downto 0); 
signal s313	: std_logic_vector(31 downto 0); 
signal s314	: std_logic_vector(31 downto 0); 
signal s315	: std_logic_vector(31 downto 0); 
signal s316	: std_logic_vector(31 downto 0); 
signal s317	: std_logic_vector(31 downto 0); 
signal s318	: std_logic_vector(31 downto 0); 
signal s319	: std_logic_vector(31 downto 0); 
signal s320	: std_logic_vector(31 downto 0); 
signal s321	: std_logic_vector(31 downto 0); 
signal s322	: std_logic_vector(31 downto 0); 
signal s323	: std_logic_vector(31 downto 0); 
signal s324	: std_logic_vector(31 downto 0); 
signal s325	: std_logic_vector(31 downto 0); 
signal s326	: std_logic_vector(31 downto 0); 
signal s327	: std_logic_vector(31 downto 0); 
signal s328	: std_logic_vector(31 downto 0); 
signal s329	: std_logic_vector(31 downto 0); 
signal s330	: std_logic_vector(31 downto 0); 
signal s331	: std_logic_vector(31 downto 0); 
signal s332	: std_logic_vector(31 downto 0); 
signal s333	: std_logic_vector(31 downto 0); 
signal s335	: std_logic_vector(31 downto 0); 
signal s336	: std_logic_vector(31 downto 0); 
signal s337	: std_logic_vector(31 downto 0); 
signal s338	: std_logic_vector(0 downto 0); 

begin 

\i\: counter
generic map ( 
	bits => 32,
	condition => 1,
	down => 0,
	increment => 2,
	steps => 1
)
port map ( 
	clk => \clk\,
	clk_en => s293,
	done => s294,
	input => s233,
	output => s299,
	reset => \reset\,
	step => s291,
	termination => s232
);

\i00\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s300,
	O0 => s185,
	reset => \reset\,
	we => s238(0)
);

\i01\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s302,
	O0 => s187,
	reset => \reset\,
	we => s240(0)
);

\i_21_add_op_s_num_22\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s33,
	O0 => s301
);

\i02\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s304,
	O0 => s189,
	reset => \reset\,
	we => s242(0)
);

\i_26_add_op_s_num_27\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s36,
	O0 => s303
);

\i10\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s306,
	O0 => s191,
	reset => \reset\,
	we => s244(0)
);

\i_31_add_op_s_num_32\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s39,
	O0 => s305
);

\i12\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s308,
	O0 => s193,
	reset => \reset\,
	we => s246(0)
);

\i_36_add_op_s_num_37\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s42,
	O0 => s307
);

\i20\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s310,
	O0 => s195,
	reset => \reset\,
	we => s248(0)
);

\i_41_add_op_s_num_42\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s45,
	O0 => s309
);

\i21\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s312,
	O0 => s197,
	reset => \reset\,
	we => s250(0)
);

\i_46_add_op_s_num_47\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s48,
	O0 => s311
);

\i22\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s314,
	O0 => s199,
	reset => \reset\,
	we => s252(0)
);

\i_51_add_op_s_num_52\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s51,
	O0 => s313
);

\H\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s52,
	O0 => s201,
	reset => \reset\,
	we => s254(0)
);

\comp_55_add_op_s_comp_62\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s53,
	I1 => s60,
	O0 => s52
);

\comp_56_add_op_s_comp_58\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s54,
	I1 => s56,
	O0 => s53
);

\i00_57_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s185,
	O0 => s54
);

\comp_59_sub_op_s_i01_61\: sub_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s57,
	I1 => s187,
	O0 => s56
);

\i01_60_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s187,
	O0 => s57
);

\comp_63_add_op_s_comp_67\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s61,
	I1 => s65,
	O0 => s60
);

\comp_64_add_op_s_i20_66\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s62,
	I1 => s195,
	O0 => s61
);

\i02_65_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s189,
	O0 => s62
);

\comp_68_add_op_s_i22_71\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s66,
	I1 => s199,
	O0 => s65
);

\i21_69_add_op_s_i21_70\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s197,
	I1 => s197,
	O0 => s66
);

\V\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s70,
	O0 => s204,
	reset => \reset\,
	we => s256(0)
);

\comp_74_add_op_s_comp_78\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s71,
	I1 => s75,
	O0 => s70
);

\comp_75_add_op_s_i02_77\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s72,
	I1 => s189,
	O0 => s71
);

\i00_76_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s185,
	O0 => s72
);

\comp_79_add_op_s_comp_87\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s76,
	I1 => s84,
	O0 => s75
);

\comp_80_add_op_s_comp_84\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s77,
	I1 => s81,
	O0 => s76
);

\comp_81_sub_op_s_i10_83\: sub_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s78,
	I1 => s191,
	O0 => s77
);

\i10_82_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s191,
	O0 => s78
);

\i12_85_add_op_s_i12_86\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s193,
	I1 => s193,
	O0 => s81
);

\comp_88_add_op_s_i22_90\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s85,
	I1 => s199,
	O0 => s84
);

\i20_89_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s195,
	O0 => s85
);

\if_lt_op_s_91\: if_lt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s201,
	I1 => s9,
	O0 => s168
);

\H_96_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s201,
	O0 => s166
);

\if_lt_op_s_97\: if_lt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s204,
	I1 => s11,
	O0 => s171
);

\V_102_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s204,
	O0 => s169
);

\O\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s92,
	O0 => s206,
	reset => \reset\,
	we => s258(0)
);

\H_105_add_op_s_V_106\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s202,
	I1 => s205,
	O0 => s92
);

\H_209\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s201,
	I1 => s166,
	O0 => s202,
	reset => \reset\,
	Sel1 => s168,
	we => s260(0)
);

\V_211\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s204,
	I1 => s169,
	O0 => s205,
	reset => \reset\,
	Sel1 => s171,
	we => s262(0)
);

\if_gt_op_s_107\: if_gt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s206,
	I1 => s13,
	O0 => s174
);

\O_213\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s206,
	I1 => s172,
	O0 => s332,
	reset => \reset\,
	Sel1 => s174,
	we => s264(0)
);

\i00_115\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s316,
	O0 => s209,
	reset => \reset\,
	we => s266(0)
);

\i_118_add_op_s_num_119\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s299,
	I1 => s106,
	O0 => s315
);

\i01_120\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s318,
	O0 => s211,
	reset => \reset\,
	we => s268(0)
);

\comp_117_add_op_s_num_123\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s108,
	O0 => s317
);

\i02_124\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s320,
	O0 => s213,
	reset => \reset\,
	we => s270(0)
);

\comp_117_add_op_s_num_127\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s110,
	O0 => s319
);

\i10_128\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s322,
	O0 => s215,
	reset => \reset\,
	we => s272(0)
);

\comp_117_add_op_s_num_131\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s112,
	O0 => s321
);

\i12_132\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s324,
	O0 => s217,
	reset => \reset\,
	we => s274(0)
);

\comp_117_add_op_s_num_135\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s114,
	O0 => s323
);

\i20_136\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s326,
	O0 => s219,
	reset => \reset\,
	we => s276(0)
);

\comp_117_add_op_s_num_139\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s116,
	O0 => s325
);

\i21_140\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s328,
	O0 => s221,
	reset => \reset\,
	we => s278(0)
);

\comp_117_add_op_s_num_143\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s118,
	O0 => s327
);

\i22_144\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s330,
	O0 => s223,
	reset => \reset\,
	we => s280(0)
);

\comp_117_add_op_s_num_147\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s315,
	I1 => s120,
	O0 => s329
);

\H_148\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s121,
	O0 => s225,
	reset => \reset\,
	we => s282(0)
);

\comp_150_add_op_s_comp_157\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s122,
	I1 => s129,
	O0 => s121
);

\comp_151_add_op_s_comp_153\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s123,
	I1 => s125,
	O0 => s122
);

\i00_152_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s209,
	O0 => s123
);

\comp_154_sub_op_s_i01_156\: sub_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s126,
	I1 => s211,
	O0 => s125
);

\i01_155_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s211,
	O0 => s126
);

\comp_158_add_op_s_comp_162\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s130,
	I1 => s134,
	O0 => s129
);

\comp_159_add_op_s_i20_161\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s131,
	I1 => s219,
	O0 => s130
);

\i02_160_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s213,
	O0 => s131
);

\comp_163_add_op_s_i22_166\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s135,
	I1 => s223,
	O0 => s134
);

\i21_164_add_op_s_i21_165\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s221,
	I1 => s221,
	O0 => s135
);

\V_167\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s139,
	O0 => s228,
	reset => \reset\,
	we => s284(0)
);

\comp_169_add_op_s_comp_173\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s140,
	I1 => s144,
	O0 => s139
);

\comp_170_add_op_s_i02_172\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s141,
	I1 => s213,
	O0 => s140
);

\i00_171_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s209,
	O0 => s141
);

\comp_174_add_op_s_comp_182\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s145,
	I1 => s153,
	O0 => s144
);

\comp_175_add_op_s_comp_179\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s146,
	I1 => s150,
	O0 => s145
);

\comp_176_sub_op_s_i10_178\: sub_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s147,
	I1 => s215,
	O0 => s146
);

\i10_177_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s215,
	O0 => s147
);

\i12_180_add_op_s_i12_181\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s217,
	I1 => s217,
	O0 => s150
);

\comp_183_add_op_s_i22_185\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s154,
	I1 => s223,
	O0 => s153
);

\i20_184_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s219,
	O0 => s154
);

\if_lt_op_s_186\: if_lt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s225,
	I1 => s24,
	O0 => s177
);

\H_191_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s225,
	O0 => s175
);

\if_lt_op_s_192\: if_lt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s228,
	I1 => s26,
	O0 => s180
);

\V_197_neg_op_s\: neg_op_s
generic map ( 
	w_in => 32,
	w_out => 32
)
port map ( 
	I0 => s228,
	O0 => s178
);

\O_198\: reg_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s161,
	O0 => s230,
	reset => \reset\,
	we => s286(0)
);

\H_200_add_op_s_V_201\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s226,
	I1 => s229,
	O0 => s161
);

\H_215\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s225,
	I1 => s175,
	O0 => s226,
	reset => \reset\,
	Sel1 => s177,
	we => s288(0)
);

\V_217\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s228,
	I1 => s178,
	O0 => s229,
	reset => \reset\,
	Sel1 => s180,
	we => s290(0)
);

\if_gt_op_s_202\: if_gt_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 1
)
port map ( 
	I0 => s230,
	I1 => s28,
	O0 => s183
);

\O_219\: reg_mux_op
generic map ( 
	initial => 0,
	w_in => 32
)
port map ( 
	clk => \clk\,
	I0 => s230,
	I1 => s181,
	O0 => s336,
	reset => \reset\,
	Sel1 => s183,
	we => s292(0)
);

\dly_225\: delay_op
generic map ( 
	bits => 32,
	delay => 7
)
port map ( 
	a => s299,
	a_delayed => s331,
	clk => \clk\,
	reset => \reset\
);

\dly_226\: delay_op
generic map ( 
	bits => 1,
	delay => 7
)
port map ( 
	a(0) => s291,
	a_delayed => s338,
	clk => \clk\,
	reset => \reset\
);

\dly_227\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s238,
	clk => \clk\,
	reset => \reset\
);

\dly_228\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s240,
	clk => \clk\,
	reset => \reset\
);

\dly_229\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s242,
	clk => \clk\,
	reset => \reset\
);

\dly_230\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s244,
	clk => \clk\,
	reset => \reset\
);

\dly_231\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s246,
	clk => \clk\,
	reset => \reset\
);

\dly_232\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s248,
	clk => \clk\,
	reset => \reset\
);

\dly_233\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s250,
	clk => \clk\,
	reset => \reset\
);

\dly_234\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s252,
	clk => \clk\,
	reset => \reset\
);

\dly_235\: delay_op
generic map ( 
	bits => 1,
	delay => 3
)
port map ( 
	a(0) => s291,
	a_delayed => s254,
	clk => \clk\,
	reset => \reset\
);

\dly_236\: delay_op
generic map ( 
	bits => 1,
	delay => 3
)
port map ( 
	a(0) => s291,
	a_delayed => s256,
	clk => \clk\,
	reset => \reset\
);

\dly_237\: delay_op
generic map ( 
	bits => 1,
	delay => 5
)
port map ( 
	a(0) => s291,
	a_delayed => s258,
	clk => \clk\,
	reset => \reset\
);

\dly_238\: delay_op
generic map ( 
	bits => 1,
	delay => 4
)
port map ( 
	a(0) => s291,
	a_delayed => s260,
	clk => \clk\,
	reset => \reset\
);

\dly_239\: delay_op
generic map ( 
	bits => 1,
	delay => 4
)
port map ( 
	a(0) => s291,
	a_delayed => s262,
	clk => \clk\,
	reset => \reset\
);

\dly_240\: delay_op
generic map ( 
	bits => 1,
	delay => 6
)
port map ( 
	a(0) => s291,
	a_delayed => s264,
	clk => \clk\,
	reset => \reset\
);

\dly_241\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s266,
	clk => \clk\,
	reset => \reset\
);

\dly_242\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s268,
	clk => \clk\,
	reset => \reset\
);

\dly_243\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s270,
	clk => \clk\,
	reset => \reset\
);

\dly_244\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s272,
	clk => \clk\,
	reset => \reset\
);

\dly_245\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s274,
	clk => \clk\,
	reset => \reset\
);

\dly_246\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s276,
	clk => \clk\,
	reset => \reset\
);

\dly_247\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s278,
	clk => \clk\,
	reset => \reset\
);

\dly_248\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s291,
	a_delayed => s280,
	clk => \clk\,
	reset => \reset\
);

\dly_249\: delay_op
generic map ( 
	bits => 1,
	delay => 3
)
port map ( 
	a(0) => s291,
	a_delayed => s282,
	clk => \clk\,
	reset => \reset\
);

\dly_250\: delay_op
generic map ( 
	bits => 1,
	delay => 3
)
port map ( 
	a(0) => s291,
	a_delayed => s284,
	clk => \clk\,
	reset => \reset\
);

\dly_251\: delay_op
generic map ( 
	bits => 1,
	delay => 5
)
port map ( 
	a(0) => s291,
	a_delayed => s286,
	clk => \clk\,
	reset => \reset\
);

\dly_252\: delay_op
generic map ( 
	bits => 1,
	delay => 4
)
port map ( 
	a(0) => s291,
	a_delayed => s288,
	clk => \clk\,
	reset => \reset\
);

\dly_253\: delay_op
generic map ( 
	bits => 1,
	delay => 4
)
port map ( 
	a(0) => s291,
	a_delayed => s290,
	clk => \clk\,
	reset => \reset\
);

\dly_254\: delay_op
generic map ( 
	bits => 1,
	delay => 6
)
port map ( 
	a(0) => s291,
	a_delayed => s292,
	clk => \clk\,
	reset => \reset\
);

\dly_255\: delay_op
generic map ( 
	bits => 1,
	delay => 9
)
port map ( 
	a(0) => s294,
	a_delayed => s295,
	clk => \clk\,
	reset => \reset\
);

\dly_256\: delay_op
generic map ( 
	bits => 32,
	delay => 7
)
port map ( 
	a => s315,
	a_delayed => s335,
	clk => \clk\,
	reset => \reset\
);

\in\: block_ram_mult_in
generic map ( 
	address_width => 7,
	data_width => 32
)
port map ( 
	address_0(6 downto 0) => s299(6 downto 0),
	data_out_0 => s300,
	address_1(6 downto 0) => s301(6 downto 0),
	data_out_1 => s302,
	address_2(6 downto 0) => s303(6 downto 0),
	data_out_2 => s304,
	address_3(6 downto 0) => s305(6 downto 0),
	data_out_3 => s306,
	address_4(6 downto 0) => s307(6 downto 0),
	data_out_4 => s308,
	address_5(6 downto 0) => s309(6 downto 0),
	data_out_5 => s310,
	address_6(6 downto 0) => s311(6 downto 0),
	data_out_6 => s312,
	address_7(6 downto 0) => s313(6 downto 0),
	data_out_7 => s314,
	address_8(6 downto 0) => s315(6 downto 0),
	data_out_8 => s316,
	address_9(6 downto 0) => s317(6 downto 0),
	data_out_9 => s318,
	address_10(6 downto 0) => s319(6 downto 0),
	data_out_10 => s320,
	address_11(6 downto 0) => s321(6 downto 0),
	data_out_11 => s322,
	address_12(6 downto 0) => s323(6 downto 0),
	data_out_12 => s324,
	address_13(6 downto 0) => s325(6 downto 0),
	data_out_13 => s326,
	address_14(6 downto 0) => s327(6 downto 0),
	data_out_14 => s328,
	address_15(6 downto 0) => s329(6 downto 0),
	data_out_15 => s330,
	clk => \clk\
);

\out\: block_ram_mult_out
generic map ( 
	address_width => 7,
	data_width => 32
)
port map ( 
	address_0(6 downto 0) => s331(6 downto 0),
	data_in_0 => s332,
	data_out_0 => s333,
	we_0 => s338(0),
	address_1(6 downto 0) => s335(6 downto 0),
	data_in_1 => s336,
	data_out_1 => s337,
	we_1 => s338(0),
	clk => \clk\
);

s33 <= conv_std_logic_vector(1, 32);
s36 <= conv_std_logic_vector(2, 32);
s39 <= conv_std_logic_vector(10, 32);
s42 <= conv_std_logic_vector(12, 32);
s45 <= conv_std_logic_vector(20, 32);
s48 <= conv_std_logic_vector(21, 32);
s51 <= conv_std_logic_vector(22, 32);
s9 <= conv_std_logic_vector(0, 32);
s11 <= conv_std_logic_vector(0, 32);
s13 <= conv_std_logic_vector(255, 32);
s172 <= conv_std_logic_vector(255, 32);
s106 <= conv_std_logic_vector(1, 32);
s108 <= conv_std_logic_vector(1, 32);
s110 <= conv_std_logic_vector(2, 32);
s112 <= conv_std_logic_vector(10, 32);
s114 <= conv_std_logic_vector(12, 32);
s116 <= conv_std_logic_vector(20, 32);
s118 <= conv_std_logic_vector(21, 32);
s120 <= conv_std_logic_vector(22, 32);
s24 <= conv_std_logic_vector(0, 32);
s26 <= conv_std_logic_vector(0, 32);
s28 <= conv_std_logic_vector(255, 32);
s181 <= conv_std_logic_vector(255, 32);
s293 <= \init\;
\done\ <= s295(0);
s232 <= conv_std_logic_vector(77, 32);
s233 <= conv_std_logic_vector(0, 32);
\out_257\ <= s333;
\out_258\ <= s337;
end behavior; 