--
-- Copyright (c) 2010 Ricardo Menotti, All Rights Reserved.
--
-- Permission to use, copy, modify, and distribute this software and its
-- documentation for NON-COMERCIAL purposes and without fee is hereby granted 
-- provided that this copyright notice appears in all copies.
--
-- RICARDO MENOTTI MAKES NO REPRESENTATIONS OR WARRANTIES ABOUT THE SUITABILITY
-- OF THE SOFTWARE, EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE, OR
-- NON-INFRINGEMENT. RICARDO MENOTTI SHALL NOT BE LIABLE FOR ANY DAMAGES
-- SUFFERED BY LICENSEE AS A RESULT OF USING, MODIFYING OR DISTRIBUTING THIS
-- SOFTWARE OR ITS DERIVATIVES.
--
-- Generated at Mon May 13 15:30:08 WEST 2013
--

-- IEEE Libraries --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity block_ram_input is
generic(
	data_width : integer := 8;
	address_width : integer := 8
);
port(
	data_in : in std_logic_vector(data_width-1 downto 0) := (others => '0');
	address : in std_logic_vector(address_width-1 downto 0);
	we: in std_logic := '0';
	oe: in std_logic := '1';
	clk : in std_logic;
	data_out : out std_logic_vector(data_width-1 downto 0));
end block_ram_input;

architecture rtl of block_ram_input is

constant mem_depth : integer := 2**address_width;
type ram_type is array (mem_depth-1 downto 0)
of std_logic_vector (data_width-1 downto 0);

signal read_a : std_logic_vector(address_width-1 downto 0);
signal RAM : ram_type := ram_type'(
	 ("0000000000000000"),	 -- 127	0
	 ("0000000000000000"),	 -- 126	0
	 ("0000000000000000"),	 -- 125	0
	 ("0000000000000000"),	 -- 124	0
	 ("0000000000000000"),	 -- 123	0
	 ("0000000000000000"),	 -- 122	0
	 ("0000000000000000"),	 -- 121	0
	 ("0000000000000000"),	 -- 120	0
	 ("0000000000000000"),	 -- 119	0
	 ("0000000000000000"),	 -- 118	0
	 ("0000000000000000"),	 -- 117	0
	 ("0000000000000000"),	 -- 116	0
	 ("0000000000000000"),	 -- 115	0
	 ("0000000000000000"),	 -- 114	0
	 ("0000000000000000"),	 -- 113	0
	 ("0000000000000000"),	 -- 112	0
	 ("0000000000000000"),	 -- 111	0
	 ("0000000000000000"),	 -- 110	0
	 ("0000000000000000"),	 -- 109	0
	 ("0000000000000000"),	 -- 108	0
	 ("0000000000000000"),	 -- 107	0
	 ("0000000000000000"),	 -- 106	0
	 ("0000000000000000"),	 -- 105	0
	 ("0000000000000000"),	 -- 104	0
	 ("0000000000000000"),	 -- 103	0
	 ("0000000000000000"),	 -- 102	0
	 ("0000000000000000"),	 -- 101	0
	 ("0000000000000000"),	 -- 100	0
	 ("0000000001100011"),	 -- 99	99
	 ("0000000000100110"),	 -- 98	38
	 ("0000000001100001"),	 -- 97	97
	 ("0000000001100000"),	 -- 96	96
	 ("0000000001011111"),	 -- 95	95
	 ("0000000001011110"),	 -- 94	94
	 ("0000000001011101"),	 -- 93	93
	 ("0000000001011100"),	 -- 92	92
	 ("0000000001100000"),	 -- 91	96
	 ("0000000001011111"),	 -- 90	95
	 ("0000000001011001"),	 -- 89	89
	 ("0000000000011100"),	 -- 88	28
	 ("0000000001010111"),	 -- 87	87
	 ("0000000001010110"),	 -- 86	86
	 ("0000000001010101"),	 -- 85	85
	 ("0000000001010100"),	 -- 84	84
	 ("0000000001010011"),	 -- 83	83
	 ("0000000001010010"),	 -- 82	82
	 ("0000000001010111"),	 -- 81	87
	 ("0000000001010100"),	 -- 80	84
	 ("0000000000011101"),	 -- 79	29
	 ("0000000000010010"),	 -- 78	18
	 ("0000000000100101"),	 -- 77	37
	 ("0000000001100000"),	 -- 76	96
	 ("0000000000110111"),	 -- 75	55
	 ("0000000000100010"),	 -- 74	34
	 ("0000000001010011"),	 -- 73	83
	 ("0000000001001000"),	 -- 72	72
	 ("0000000001000100"),	 -- 71	68
	 ("0000000000110101"),	 -- 70	53
	 ("0000000001000101"),	 -- 69	69
	 ("0000000001000100"),	 -- 68	68
	 ("0000000001000011"),	 -- 67	67
	 ("0000000001000000"),	 -- 66	64
	 ("0000000001000001"),	 -- 65	65
	 ("0000000001000000"),	 -- 64	64
	 ("0000000001000010"),	 -- 63	66
	 ("0000000000111110"),	 -- 62	62
	 ("0000000001000101"),	 -- 61	69
	 ("0000000000111100"),	 -- 60	60
	 ("0000000000011101"),	 -- 59	29
	 ("0000000000010010"),	 -- 58	18
	 ("0000000000100101"),	 -- 57	37
	 ("0000000001100000"),	 -- 56	96
	 ("0000000000101101"),	 -- 55	45
	 ("0000000000100010"),	 -- 54	34
	 ("0000000001010011"),	 -- 53	83
	 ("0000000001010010"),	 -- 52	82
	 ("0000000000111100"),	 -- 51	60
	 ("0000000000110100"),	 -- 50	52
	 ("0000000001011001"),	 -- 49	89
	 ("0000000000110000"),	 -- 48	48
	 ("0000000000101111"),	 -- 47	47
	 ("0000000000101110"),	 -- 46	46
	 ("0000000000101101"),	 -- 45	45
	 ("0000000000101100"),	 -- 44	44
	 ("0000000001001001"),	 -- 43	73
	 ("0000000000101010"),	 -- 42	42
	 ("0000000000101001"),	 -- 41	41
	 ("0000000000101000"),	 -- 40	40
	 ("0000000000011101"),	 -- 39	29
	 ("0000000000010010"),	 -- 38	18
	 ("0000000001100001"),	 -- 37	97
	 ("0000000001100000"),	 -- 36	96
	 ("0000000000101101"),	 -- 35	45
	 ("0000000000100010"),	 -- 34	34
	 ("0000000001010011"),	 -- 33	83
	 ("0000000001001000"),	 -- 32	72
	 ("0000000000001100"),	 -- 31	12
	 ("0000000000110110"),	 -- 30	54
	 ("0000000000011101"),	 -- 29	29
	 ("0000000000011100"),	 -- 28	28
	 ("0000000000011011"),	 -- 27	27
	 ("0000000000011010"),	 -- 26	26
	 ("0000000000011001"),	 -- 25	25
	 ("0000000000010100"),	 -- 24	20
	 ("0000000000010111"),	 -- 23	23
	 ("0000000001010010"),	 -- 22	82
	 ("0000000000010111"),	 -- 21	23
	 ("0000000000010100"),	 -- 20	20
	 ("0000000000100111"),	 -- 19	39
	 ("0000000000010010"),	 -- 18	18
	 ("0000000000010001"),	 -- 17	17
	 ("0000000000010000"),	 -- 16	16
	 ("0000000000001111"),	 -- 15	15
	 ("0000000000001110"),	 -- 14	14
	 ("0000000000001101"),	 -- 13	13
	 ("0000000001001000"),	 -- 12	72
	 ("0000000000001110"),	 -- 11	14
	 ("0000000000001110"),	 -- 10	14
	 ("0000000000011101"),	 -- 9	29
	 ("0000000000010010"),	 -- 8	18
	 ("0000000001000011"),	 -- 7	67
	 ("0000000001100000"),	 -- 6	96
	 ("0000000000101101"),	 -- 5	45
	 ("0000000000100010"),	 -- 4	34
	 ("0000000001010011"),	 -- 3	83
	 ("0000000000111110"),	 -- 2	62
	 ("0000000001000001"),	 -- 1	65
	 ("0000000000110010"));	 -- 0	50

begin
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we = '1') then
        RAM(conv_integer(address)) <= data_in;
        data_out <= RAM(conv_integer(read_a));
      elsif (oe = '1') then
        data_out <= RAM(conv_integer(read_a));
      end if;
      read_a <= address;
    end if;
  end process;
end rtl;
