--
-- Copyright (c) 2010 Ricardo Menotti, All Rights Reserved.
--
-- Permission to use, copy, modify, and distribute this software and its
-- documentation for NON-COMERCIAL purposes and without fee is hereby granted 
-- provided that this copyright notice appears in all copies.
--
-- RICARDO MENOTTI MAKES NO REPRESENTATIONS OR WARRANTIES ABOUT THE SUITABILITY
-- OF THE SOFTWARE, EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE, OR
-- NON-INFRINGEMENT. RICARDO MENOTTI SHALL NOT BE LIABLE FOR ANY DAMAGES
-- SUFFERED BY LICENSEE AS A RESULT OF USING, MODIFYING OR DISTRIBUTING THIS
-- SOFTWARE OR ITS DERIVATIVES.
--
-- Generated at Tue Oct 25 21:42:50 BRST 2011
--

-- IEEE Libraries --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity block_ram_dct_io_ptr is
generic(
	data_width : integer := 8;
	address_width : integer := 8
);
port(
	data_in : in std_logic_vector(data_width-1 downto 0) := (others => '0');
	address : in std_logic_vector(address_width-1 downto 0);
	we: in std_logic := '0';
	oe: in std_logic := '1';
	clk : in std_logic;
	data_out : out std_logic_vector(data_width-1 downto 0));
end block_ram_dct_io_ptr;

architecture rtl of block_ram_dct_io_ptr is

constant mem_depth : integer := 2**address_width;
type ram_type is array (mem_depth-1 downto 0)
of std_logic_vector (data_width-1 downto 0);

signal read_a : std_logic_vector(address_width-1 downto 0);
signal RAM : ram_type := ram_type'(
	 ("00000000000000000000000000000000"),	 -- 1023	0
	 ("00000000000000000000000000000000"),	 -- 1022	0
	 ("00000000000000000000000000000000"),	 -- 1021	0
	 ("00000000000000000000000000000000"),	 -- 1020	0
	 ("00000000000000000000000000000000"),	 -- 1019	0
	 ("00000000000000000000000000000000"),	 -- 1018	0
	 ("00000000000000000000000000000000"),	 -- 1017	0
	 ("00000000000000000000000000000000"),	 -- 1016	0
	 ("00000000000000000000000000000000"),	 -- 1015	0
	 ("00000000000000000000000000000000"),	 -- 1014	0
	 ("00000000000000000000000000000000"),	 -- 1013	0
	 ("00000000000000000000000000000000"),	 -- 1012	0
	 ("00000000000000000000000000000000"),	 -- 1011	0
	 ("00000000000000000000000000000000"),	 -- 1010	0
	 ("00000000000000000000000000000000"),	 -- 1009	0
	 ("00000000000000000000000000000000"),	 -- 1008	0
	 ("00000000000000000000000000000000"),	 -- 1007	0
	 ("00000000000000000000000000000000"),	 -- 1006	0
	 ("00000000000000000000000000000000"),	 -- 1005	0
	 ("00000000000000000000000000000000"),	 -- 1004	0
	 ("00000000000000000000000000000000"),	 -- 1003	0
	 ("00000000000000000000000000000000"),	 -- 1002	0
	 ("00000000000000000000000000000000"),	 -- 1001	0
	 ("00000000000000000000000000000000"),	 -- 1000	0
	 ("00000000000000000000000000000000"),	 -- 999	0
	 ("00000000000000000000000000000000"),	 -- 998	0
	 ("00000000000000000000000000000000"),	 -- 997	0
	 ("00000000000000000000000000000000"),	 -- 996	0
	 ("00000000000000000000000000000000"),	 -- 995	0
	 ("00000000000000000000000000000000"),	 -- 994	0
	 ("00000000000000000000000000000000"),	 -- 993	0
	 ("00000000000000000000000000000000"),	 -- 992	0
	 ("00000000000000000000000000000000"),	 -- 991	0
	 ("00000000000000000000000000000000"),	 -- 990	0
	 ("00000000000000000000000000000000"),	 -- 989	0
	 ("00000000000000000000000000000000"),	 -- 988	0
	 ("00000000000000000000000000000000"),	 -- 987	0
	 ("00000000000000000000000000000000"),	 -- 986	0
	 ("00000000000000000000000000000000"),	 -- 985	0
	 ("00000000000000000000000000000000"),	 -- 984	0
	 ("00000000000000000000000000000000"),	 -- 983	0
	 ("00000000000000000000000000000000"),	 -- 982	0
	 ("00000000000000000000000000000000"),	 -- 981	0
	 ("00000000000000000000000000000000"),	 -- 980	0
	 ("00000000000000000000000000000000"),	 -- 979	0
	 ("00000000000000000000000000000000"),	 -- 978	0
	 ("00000000000000000000000000000000"),	 -- 977	0
	 ("00000000000000000000000000000000"),	 -- 976	0
	 ("00000000000000000000000000000000"),	 -- 975	0
	 ("00000000000000000000000000000000"),	 -- 974	0
	 ("00000000000000000000000000000000"),	 -- 973	0
	 ("00000000000000000000000000000000"),	 -- 972	0
	 ("00000000000000000000000000000000"),	 -- 971	0
	 ("00000000000000000000000000000000"),	 -- 970	0
	 ("00000000000000000000000000000000"),	 -- 969	0
	 ("00000000000000000000000000000000"),	 -- 968	0
	 ("00000000000000000000000000000000"),	 -- 967	0
	 ("00000000000000000000000000000000"),	 -- 966	0
	 ("00000000000000000000000000000000"),	 -- 965	0
	 ("00000000000000000000000000000000"),	 -- 964	0
	 ("00000000000000000000000000000000"),	 -- 963	0
	 ("00000000000000000000000000000000"),	 -- 962	0
	 ("00000000000000000000000000000000"),	 -- 961	0
	 ("00000000000000000000000000000000"),	 -- 960	0
	 ("00000000000000000000000000000000"),	 -- 959	0
	 ("00000000000000000000000000000000"),	 -- 958	0
	 ("00000000000000000000000000000000"),	 -- 957	0
	 ("00000000000000000000000000000000"),	 -- 956	0
	 ("00000000000000000000000000000000"),	 -- 955	0
	 ("00000000000000000000000000000000"),	 -- 954	0
	 ("00000000000000000000000000000000"),	 -- 953	0
	 ("00000000000000000000000000000000"),	 -- 952	0
	 ("00000000000000000000000000000000"),	 -- 951	0
	 ("00000000000000000000000000000000"),	 -- 950	0
	 ("00000000000000000000000000000000"),	 -- 949	0
	 ("00000000000000000000000000000000"),	 -- 948	0
	 ("00000000000000000000000000000000"),	 -- 947	0
	 ("00000000000000000000000000000000"),	 -- 946	0
	 ("00000000000000000000000000000000"),	 -- 945	0
	 ("00000000000000000000000000000000"),	 -- 944	0
	 ("00000000000000000000000000000000"),	 -- 943	0
	 ("00000000000000000000000000000000"),	 -- 942	0
	 ("00000000000000000000000000000000"),	 -- 941	0
	 ("00000000000000000000000000000000"),	 -- 940	0
	 ("00000000000000000000000000000000"),	 -- 939	0
	 ("00000000000000000000000000000000"),	 -- 938	0
	 ("00000000000000000000000000000000"),	 -- 937	0
	 ("00000000000000000000000000000000"),	 -- 936	0
	 ("00000000000000000000000000000000"),	 -- 935	0
	 ("00000000000000000000000000000000"),	 -- 934	0
	 ("00000000000000000000000000000000"),	 -- 933	0
	 ("00000000000000000000000000000000"),	 -- 932	0
	 ("00000000000000000000000000000000"),	 -- 931	0
	 ("00000000000000000000000000000000"),	 -- 930	0
	 ("00000000000000000000000000000000"),	 -- 929	0
	 ("00000000000000000000000000000000"),	 -- 928	0
	 ("00000000000000000000000000000000"),	 -- 927	0
	 ("00000000000000000000000000000000"),	 -- 926	0
	 ("00000000000000000000000000000000"),	 -- 925	0
	 ("00000000000000000000000000000000"),	 -- 924	0
	 ("00000000000000000000000000000000"),	 -- 923	0
	 ("00000000000000000000000000000000"),	 -- 922	0
	 ("00000000000000000000000000000000"),	 -- 921	0
	 ("00000000000000000000000000000000"),	 -- 920	0
	 ("00000000000000000000000000000000"),	 -- 919	0
	 ("00000000000000000000000000000000"),	 -- 918	0
	 ("00000000000000000000000000000000"),	 -- 917	0
	 ("00000000000000000000000000000000"),	 -- 916	0
	 ("00000000000000000000000000000000"),	 -- 915	0
	 ("00000000000000000000000000000000"),	 -- 914	0
	 ("00000000000000000000000000000000"),	 -- 913	0
	 ("00000000000000000000000000000000"),	 -- 912	0
	 ("00000000000000000000000000000000"),	 -- 911	0
	 ("00000000000000000000000000000000"),	 -- 910	0
	 ("00000000000000000000000000000000"),	 -- 909	0
	 ("00000000000000000000000000000000"),	 -- 908	0
	 ("00000000000000000000000000000000"),	 -- 907	0
	 ("00000000000000000000000000000000"),	 -- 906	0
	 ("00000000000000000000000000000000"),	 -- 905	0
	 ("00000000000000000000000000000000"),	 -- 904	0
	 ("00000000000000000000000000000000"),	 -- 903	0
	 ("00000000000000000000000000000000"),	 -- 902	0
	 ("00000000000000000000000000000000"),	 -- 901	0
	 ("00000000000000000000000000000000"),	 -- 900	0
	 ("00000000000000000000000000000000"),	 -- 899	0
	 ("00000000000000000000000000000000"),	 -- 898	0
	 ("00000000000000000000000000000000"),	 -- 897	0
	 ("00000000000000000000000000000000"),	 -- 896	0
	 ("00000000000000000000000000000000"),	 -- 895	0
	 ("00000000000000000000000000000000"),	 -- 894	0
	 ("00000000000000000000000000000000"),	 -- 893	0
	 ("00000000000000000000000000000000"),	 -- 892	0
	 ("00000000000000000000000000000000"),	 -- 891	0
	 ("00000000000000000000000000000000"),	 -- 890	0
	 ("00000000000000000000000000000000"),	 -- 889	0
	 ("00000000000000000000000000000000"),	 -- 888	0
	 ("00000000000000000000000000000000"),	 -- 887	0
	 ("00000000000000000000000000000000"),	 -- 886	0
	 ("00000000000000000000000000000000"),	 -- 885	0
	 ("00000000000000000000000000000000"),	 -- 884	0
	 ("00000000000000000000000000000000"),	 -- 883	0
	 ("00000000000000000000000000000000"),	 -- 882	0
	 ("00000000000000000000000000000000"),	 -- 881	0
	 ("00000000000000000000000000000000"),	 -- 880	0
	 ("00000000000000000000000000000000"),	 -- 879	0
	 ("00000000000000000000000000000000"),	 -- 878	0
	 ("00000000000000000000000000000000"),	 -- 877	0
	 ("00000000000000000000000000000000"),	 -- 876	0
	 ("00000000000000000000000000000000"),	 -- 875	0
	 ("00000000000000000000000000000000"),	 -- 874	0
	 ("00000000000000000000000000000000"),	 -- 873	0
	 ("00000000000000000000000000000000"),	 -- 872	0
	 ("00000000000000000000000000000000"),	 -- 871	0
	 ("00000000000000000000000000000000"),	 -- 870	0
	 ("00000000000000000000000000000000"),	 -- 869	0
	 ("00000000000000000000000000000000"),	 -- 868	0
	 ("00000000000000000000000000000000"),	 -- 867	0
	 ("00000000000000000000000000000000"),	 -- 866	0
	 ("00000000000000000000000000000000"),	 -- 865	0
	 ("00000000000000000000000000000000"),	 -- 864	0
	 ("00000000000000000000000000000000"),	 -- 863	0
	 ("00000000000000000000000000000000"),	 -- 862	0
	 ("00000000000000000000000000000000"),	 -- 861	0
	 ("00000000000000000000000000000000"),	 -- 860	0
	 ("00000000000000000000000000000000"),	 -- 859	0
	 ("00000000000000000000000000000000"),	 -- 858	0
	 ("00000000000000000000000000000000"),	 -- 857	0
	 ("00000000000000000000000000000000"),	 -- 856	0
	 ("00000000000000000000000000000000"),	 -- 855	0
	 ("00000000000000000000000000000000"),	 -- 854	0
	 ("00000000000000000000000000000000"),	 -- 853	0
	 ("00000000000000000000000000000000"),	 -- 852	0
	 ("00000000000000000000000000000000"),	 -- 851	0
	 ("00000000000000000000000000000000"),	 -- 850	0
	 ("00000000000000000000000000000000"),	 -- 849	0
	 ("00000000000000000000000000000000"),	 -- 848	0
	 ("00000000000000000000000000000000"),	 -- 847	0
	 ("00000000000000000000000000000000"),	 -- 846	0
	 ("00000000000000000000000000000000"),	 -- 845	0
	 ("00000000000000000000000000000000"),	 -- 844	0
	 ("00000000000000000000000000000000"),	 -- 843	0
	 ("00000000000000000000000000000000"),	 -- 842	0
	 ("00000000000000000000000000000000"),	 -- 841	0
	 ("00000000000000000000000000000000"),	 -- 840	0
	 ("00000000000000000000000000000000"),	 -- 839	0
	 ("00000000000000000000000000000000"),	 -- 838	0
	 ("00000000000000000000000000000000"),	 -- 837	0
	 ("00000000000000000000000000000000"),	 -- 836	0
	 ("00000000000000000000000000000000"),	 -- 835	0
	 ("00000000000000000000000000000000"),	 -- 834	0
	 ("00000000000000000000000000000000"),	 -- 833	0
	 ("00000000000000000000000000000000"),	 -- 832	0
	 ("00000000000000000000000000000000"),	 -- 831	0
	 ("00000000000000000000000000000000"),	 -- 830	0
	 ("00000000000000000000000000000000"),	 -- 829	0
	 ("00000000000000000000000000000000"),	 -- 828	0
	 ("00000000000000000000000000000000"),	 -- 827	0
	 ("00000000000000000000000000000000"),	 -- 826	0
	 ("00000000000000000000000000000000"),	 -- 825	0
	 ("00000000000000000000000000000000"),	 -- 824	0
	 ("00000000000000000000000000000000"),	 -- 823	0
	 ("00000000000000000000000000000000"),	 -- 822	0
	 ("00000000000000000000000000000000"),	 -- 821	0
	 ("00000000000000000000000000000000"),	 -- 820	0
	 ("00000000000000000000000000000000"),	 -- 819	0
	 ("00000000000000000000000000000000"),	 -- 818	0
	 ("00000000000000000000000000000000"),	 -- 817	0
	 ("00000000000000000000000000000000"),	 -- 816	0
	 ("00000000000000000000000000000000"),	 -- 815	0
	 ("00000000000000000000000000000000"),	 -- 814	0
	 ("00000000000000000000000000000000"),	 -- 813	0
	 ("00000000000000000000000000000000"),	 -- 812	0
	 ("00000000000000000000000000000000"),	 -- 811	0
	 ("00000000000000000000000000000000"),	 -- 810	0
	 ("00000000000000000000000000000000"),	 -- 809	0
	 ("00000000000000000000000000000000"),	 -- 808	0
	 ("00000000000000000000000000000000"),	 -- 807	0
	 ("00000000000000000000000000000000"),	 -- 806	0
	 ("00000000000000000000000000000000"),	 -- 805	0
	 ("00000000000000000000000000000000"),	 -- 804	0
	 ("00000000000000000000000000000000"),	 -- 803	0
	 ("00000000000000000000000000000000"),	 -- 802	0
	 ("00000000000000000000000000000000"),	 -- 801	0
	 ("00000000000000000000000000000000"),	 -- 800	0
	 ("00000000000000000000000000000000"),	 -- 799	0
	 ("00000000000000000000000000000000"),	 -- 798	0
	 ("00000000000000000000000000000000"),	 -- 797	0
	 ("00000000000000000000000000000000"),	 -- 796	0
	 ("00000000000000000000000000000000"),	 -- 795	0
	 ("00000000000000000000000000000000"),	 -- 794	0
	 ("00000000000000000000000000000000"),	 -- 793	0
	 ("00000000000000000000000000000000"),	 -- 792	0
	 ("00000000000000000000000000000000"),	 -- 791	0
	 ("00000000000000000000000000000000"),	 -- 790	0
	 ("00000000000000000000000000000000"),	 -- 789	0
	 ("00000000000000000000000000000000"),	 -- 788	0
	 ("00000000000000000000000000000000"),	 -- 787	0
	 ("00000000000000000000000000000000"),	 -- 786	0
	 ("00000000000000000000000000000000"),	 -- 785	0
	 ("00000000000000000000000000000000"),	 -- 784	0
	 ("00000000000000000000000000000000"),	 -- 783	0
	 ("00000000000000000000000000000000"),	 -- 782	0
	 ("00000000000000000000000000000000"),	 -- 781	0
	 ("00000000000000000000000000000000"),	 -- 780	0
	 ("00000000000000000000000000000000"),	 -- 779	0
	 ("00000000000000000000000000000000"),	 -- 778	0
	 ("00000000000000000000000000000000"),	 -- 777	0
	 ("00000000000000000000000000000000"),	 -- 776	0
	 ("00000000000000000000000000000000"),	 -- 775	0
	 ("00000000000000000000000000000000"),	 -- 774	0
	 ("00000000000000000000000000000000"),	 -- 773	0
	 ("00000000000000000000000000000000"),	 -- 772	0
	 ("00000000000000000000000000000000"),	 -- 771	0
	 ("00000000000000000000000000000000"),	 -- 770	0
	 ("00000000000000000000000000000000"),	 -- 769	0
	 ("00000000000000000000000000000000"),	 -- 768	0
	 ("00000000000000000000000000000000"),	 -- 767	0
	 ("00000000000000000000000000000000"),	 -- 766	0
	 ("00000000000000000000000000000000"),	 -- 765	0
	 ("00000000000000000000000000000000"),	 -- 764	0
	 ("00000000000000000000000000000000"),	 -- 763	0
	 ("00000000000000000000000000000000"),	 -- 762	0
	 ("00000000000000000000000000000000"),	 -- 761	0
	 ("00000000000000000000000000000000"),	 -- 760	0
	 ("00000000000000000000000000000000"),	 -- 759	0
	 ("00000000000000000000000000000000"),	 -- 758	0
	 ("00000000000000000000000000000000"),	 -- 757	0
	 ("00000000000000000000000000000000"),	 -- 756	0
	 ("00000000000000000000000000000000"),	 -- 755	0
	 ("00000000000000000000000000000000"),	 -- 754	0
	 ("00000000000000000000000000000000"),	 -- 753	0
	 ("00000000000000000000000000000000"),	 -- 752	0
	 ("00000000000000000000000000000000"),	 -- 751	0
	 ("00000000000000000000000000000000"),	 -- 750	0
	 ("00000000000000000000000000000000"),	 -- 749	0
	 ("00000000000000000000000000000000"),	 -- 748	0
	 ("00000000000000000000000000000000"),	 -- 747	0
	 ("00000000000000000000000000000000"),	 -- 746	0
	 ("00000000000000000000000000000000"),	 -- 745	0
	 ("00000000000000000000000000000000"),	 -- 744	0
	 ("00000000000000000000000000000000"),	 -- 743	0
	 ("00000000000000000000000000000000"),	 -- 742	0
	 ("00000000000000000000000000000000"),	 -- 741	0
	 ("00000000000000000000000000000000"),	 -- 740	0
	 ("00000000000000000000000000000000"),	 -- 739	0
	 ("00000000000000000000000000000000"),	 -- 738	0
	 ("00000000000000000000000000000000"),	 -- 737	0
	 ("00000000000000000000000000000000"),	 -- 736	0
	 ("00000000000000000000000000000000"),	 -- 735	0
	 ("00000000000000000000000000000000"),	 -- 734	0
	 ("00000000000000000000000000000000"),	 -- 733	0
	 ("00000000000000000000000000000000"),	 -- 732	0
	 ("00000000000000000000000000000000"),	 -- 731	0
	 ("00000000000000000000000000000000"),	 -- 730	0
	 ("00000000000000000000000000000000"),	 -- 729	0
	 ("00000000000000000000000000000000"),	 -- 728	0
	 ("00000000000000000000000000000000"),	 -- 727	0
	 ("00000000000000000000000000000000"),	 -- 726	0
	 ("00000000000000000000000000000000"),	 -- 725	0
	 ("00000000000000000000000000000000"),	 -- 724	0
	 ("00000000000000000000000000000000"),	 -- 723	0
	 ("00000000000000000000000000000000"),	 -- 722	0
	 ("00000000000000000000000000000000"),	 -- 721	0
	 ("00000000000000000000000000000000"),	 -- 720	0
	 ("00000000000000000000000000000000"),	 -- 719	0
	 ("00000000000000000000000000000000"),	 -- 718	0
	 ("00000000000000000000000000000000"),	 -- 717	0
	 ("00000000000000000000000000000000"),	 -- 716	0
	 ("00000000000000000000000000000000"),	 -- 715	0
	 ("00000000000000000000000000000000"),	 -- 714	0
	 ("00000000000000000000000000000000"),	 -- 713	0
	 ("00000000000000000000000000000000"),	 -- 712	0
	 ("00000000000000000000000000000000"),	 -- 711	0
	 ("00000000000000000000000000000000"),	 -- 710	0
	 ("00000000000000000000000000000000"),	 -- 709	0
	 ("00000000000000000000000000000000"),	 -- 708	0
	 ("00000000000000000000000000000000"),	 -- 707	0
	 ("00000000000000000000000000000000"),	 -- 706	0
	 ("00000000000000000000000000000000"),	 -- 705	0
	 ("00000000000000000000000000000000"),	 -- 704	0
	 ("00000000000000000000000000000000"),	 -- 703	0
	 ("00000000000000000000000000000000"),	 -- 702	0
	 ("00000000000000000000000000000000"),	 -- 701	0
	 ("00000000000000000000000000000000"),	 -- 700	0
	 ("00000000000000000000000000000000"),	 -- 699	0
	 ("00000000000000000000000000000000"),	 -- 698	0
	 ("00000000000000000000000000000000"),	 -- 697	0
	 ("00000000000000000000000000000000"),	 -- 696	0
	 ("00000000000000000000000000000000"),	 -- 695	0
	 ("00000000000000000000000000000000"),	 -- 694	0
	 ("00000000000000000000000000000000"),	 -- 693	0
	 ("00000000000000000000000000000000"),	 -- 692	0
	 ("00000000000000000000000000000000"),	 -- 691	0
	 ("00000000000000000000000000000000"),	 -- 690	0
	 ("00000000000000000000000000000000"),	 -- 689	0
	 ("00000000000000000000000000000000"),	 -- 688	0
	 ("00000000000000000000000000000000"),	 -- 687	0
	 ("00000000000000000000000000000000"),	 -- 686	0
	 ("00000000000000000000000000000000"),	 -- 685	0
	 ("00000000000000000000000000000000"),	 -- 684	0
	 ("00000000000000000000000000000000"),	 -- 683	0
	 ("00000000000000000000000000000000"),	 -- 682	0
	 ("00000000000000000000000000000000"),	 -- 681	0
	 ("00000000000000000000000000000000"),	 -- 680	0
	 ("00000000000000000000000000000000"),	 -- 679	0
	 ("00000000000000000000000000000000"),	 -- 678	0
	 ("00000000000000000000000000000000"),	 -- 677	0
	 ("00000000000000000000000000000000"),	 -- 676	0
	 ("00000000000000000000000000000000"),	 -- 675	0
	 ("00000000000000000000000000000000"),	 -- 674	0
	 ("00000000000000000000000000000000"),	 -- 673	0
	 ("00000000000000000000000000000000"),	 -- 672	0
	 ("00000000000000000000000000000000"),	 -- 671	0
	 ("00000000000000000000000000000000"),	 -- 670	0
	 ("00000000000000000000000000000000"),	 -- 669	0
	 ("00000000000000000000000000000000"),	 -- 668	0
	 ("00000000000000000000000000000000"),	 -- 667	0
	 ("00000000000000000000000000000000"),	 -- 666	0
	 ("00000000000000000000000000000000"),	 -- 665	0
	 ("00000000000000000000000000000000"),	 -- 664	0
	 ("00000000000000000000000000000000"),	 -- 663	0
	 ("00000000000000000000000000000000"),	 -- 662	0
	 ("00000000000000000000000000000000"),	 -- 661	0
	 ("00000000000000000000000000000000"),	 -- 660	0
	 ("00000000000000000000000000000000"),	 -- 659	0
	 ("00000000000000000000000000000000"),	 -- 658	0
	 ("00000000000000000000000000000000"),	 -- 657	0
	 ("00000000000000000000000000000000"),	 -- 656	0
	 ("00000000000000000000000000000000"),	 -- 655	0
	 ("00000000000000000000000000000000"),	 -- 654	0
	 ("00000000000000000000000000000000"),	 -- 653	0
	 ("00000000000000000000000000000000"),	 -- 652	0
	 ("00000000000000000000000000000000"),	 -- 651	0
	 ("00000000000000000000000000000000"),	 -- 650	0
	 ("00000000000000000000000000000000"),	 -- 649	0
	 ("00000000000000000000000000000000"),	 -- 648	0
	 ("00000000000000000000000000000000"),	 -- 647	0
	 ("00000000000000000000000000000000"),	 -- 646	0
	 ("00000000000000000000000000000000"),	 -- 645	0
	 ("00000000000000000000000000000000"),	 -- 644	0
	 ("00000000000000000000000000000000"),	 -- 643	0
	 ("00000000000000000000000000000000"),	 -- 642	0
	 ("00000000000000000000000000000000"),	 -- 641	0
	 ("00000000000000000000000000000000"),	 -- 640	0
	 ("00000000000000000000000110010111"),	 -- 639	407
	 ("11111111111111111111101000011100"),	 -- 638	-1508
	 ("00000000000000000000000110010101"),	 -- 637	405
	 ("00000000000000000000000110010100"),	 -- 636	404
	 ("11111111111111111111101000100010"),	 -- 635	-1502
	 ("00000000000000000000000110010010"),	 -- 634	402
	 ("00000000000000000000000110010001"),	 -- 633	401
	 ("11111111111111111111101000101000"),	 -- 632	-1496
	 ("00000000000000000000000110001111"),	 -- 631	399
	 ("00000000000000000000000110001110"),	 -- 630	398
	 ("11111111111111111111101000101110"),	 -- 629	-1490
	 ("00000000000000000000000110001100"),	 -- 628	396
	 ("00000000000000000000000110001011"),	 -- 627	395
	 ("11111111111111111111101000110100"),	 -- 626	-1484
	 ("00000000000000000000000110001001"),	 -- 625	393
	 ("00000000000000000000000110001000"),	 -- 624	392
	 ("11111111111111111111101000111010"),	 -- 623	-1478
	 ("00000000000000000000000110000110"),	 -- 622	390
	 ("00000000000000000000000110000101"),	 -- 621	389
	 ("11111111111111111111101001000000"),	 -- 620	-1472
	 ("00000000000000000000000110000011"),	 -- 619	387
	 ("00000000000000000000000110000010"),	 -- 618	386
	 ("11111111111111111111101001000110"),	 -- 617	-1466
	 ("00000000000000000000000110000000"),	 -- 616	384
	 ("00000000000000000000000101111111"),	 -- 615	383
	 ("11111111111111111111101001001100"),	 -- 614	-1460
	 ("00000000000000000000000101111101"),	 -- 613	381
	 ("00000000000000000000000101111100"),	 -- 612	380
	 ("11111111111111111111101001010010"),	 -- 611	-1454
	 ("00000000000000000000000101111010"),	 -- 610	378
	 ("00000000000000000000000101111001"),	 -- 609	377
	 ("11111111111111111111101001011000"),	 -- 608	-1448
	 ("00000000000000000000000101110111"),	 -- 607	375
	 ("00000000000000000000000101110110"),	 -- 606	374
	 ("11111111111111111111101001011110"),	 -- 605	-1442
	 ("00000000000000000000000101110100"),	 -- 604	372
	 ("00000000000000000000000101110011"),	 -- 603	371
	 ("11111111111111111111101001100100"),	 -- 602	-1436
	 ("00000000000000000000000101110001"),	 -- 601	369
	 ("00000000000000000000000101110000"),	 -- 600	368
	 ("11111111111111111111101001101010"),	 -- 599	-1430
	 ("00000000000000000000000101101110"),	 -- 598	366
	 ("00000000000000000000000101101101"),	 -- 597	365
	 ("11111111111111111111101001110000"),	 -- 596	-1424
	 ("00000000000000000000000101101011"),	 -- 595	363
	 ("00000000000000000000000101101010"),	 -- 594	362
	 ("11111111111111111111101001110110"),	 -- 593	-1418
	 ("00000000000000000000000101101000"),	 -- 592	360
	 ("00000000000000000000000101100111"),	 -- 591	359
	 ("11111111111111111111101001111100"),	 -- 590	-1412
	 ("00000000000000000000000101100101"),	 -- 589	357
	 ("00000000000000000000000101100100"),	 -- 588	356
	 ("11111111111111111111101010000010"),	 -- 587	-1406
	 ("00000000000000000000000101100010"),	 -- 586	354
	 ("00000000000000000000000101100001"),	 -- 585	353
	 ("11111111111111111111101010001000"),	 -- 584	-1400
	 ("00000000000000000000000101011111"),	 -- 583	351
	 ("00000000000000000000000101011110"),	 -- 582	350
	 ("11111111111111111111101010001110"),	 -- 581	-1394
	 ("00000000000000000000000101011100"),	 -- 580	348
	 ("00000000000000000000000101011011"),	 -- 579	347
	 ("11111111111111111111101010010100"),	 -- 578	-1388
	 ("00000000000000000000000101011001"),	 -- 577	345
	 ("00000000000000000000000101011000"),	 -- 576	344
	 ("11111111111111111111101010011010"),	 -- 575	-1382
	 ("00000000000000000000000101010110"),	 -- 574	342
	 ("00000000000000000000000101010101"),	 -- 573	341
	 ("11111111111111111111101010100000"),	 -- 572	-1376
	 ("00000000000000000000000101010011"),	 -- 571	339
	 ("00000000000000000000000101010010"),	 -- 570	338
	 ("11111111111111111111101010100110"),	 -- 569	-1370
	 ("00000000000000000000000101010000"),	 -- 568	336
	 ("00000000000000000000000101001111"),	 -- 567	335
	 ("11111111111111111111101010101100"),	 -- 566	-1364
	 ("00000000000000000000000101001101"),	 -- 565	333
	 ("00000000000000000000000101001100"),	 -- 564	332
	 ("11111111111111111111101010110010"),	 -- 563	-1358
	 ("00000000000000000000000101001010"),	 -- 562	330
	 ("00000000000000000000000101001001"),	 -- 561	329
	 ("11111111111111111111101010111000"),	 -- 560	-1352
	 ("00000000000000000000000101000111"),	 -- 559	327
	 ("00000000000000000000000101000110"),	 -- 558	326
	 ("11111111111111111111101010111110"),	 -- 557	-1346
	 ("00000000000000000000000101000100"),	 -- 556	324
	 ("00000000000000000000000101000011"),	 -- 555	323
	 ("11111111111111111111101011000100"),	 -- 554	-1340
	 ("00000000000000000000000101000001"),	 -- 553	321
	 ("00000000000000000000000101000000"),	 -- 552	320
	 ("11111111111111111111101011001010"),	 -- 551	-1334
	 ("00000000000000000000000100111110"),	 -- 550	318
	 ("00000000000000000000000100111101"),	 -- 549	317
	 ("11111111111111111111101011010000"),	 -- 548	-1328
	 ("00000000000000000000000100111011"),	 -- 547	315
	 ("00000000000000000000000100111010"),	 -- 546	314
	 ("11111111111111111111101011010110"),	 -- 545	-1322
	 ("00000000000000000000000100111000"),	 -- 544	312
	 ("00000000000000000000000100110111"),	 -- 543	311
	 ("11111111111111111111101011011100"),	 -- 542	-1316
	 ("00000000000000000000000100110101"),	 -- 541	309
	 ("00000000000000000000000100110100"),	 -- 540	308
	 ("11111111111111111111101011100010"),	 -- 539	-1310
	 ("00000000000000000000000100110010"),	 -- 538	306
	 ("00000000000000000000000100110001"),	 -- 537	305
	 ("11111111111111111111101011101000"),	 -- 536	-1304
	 ("00000000000000000000000100101111"),	 -- 535	303
	 ("00000000000000000000000100101110"),	 -- 534	302
	 ("11111111111111111111101011101110"),	 -- 533	-1298
	 ("00000000000000000000000100101100"),	 -- 532	300
	 ("00000000000000000000000100101011"),	 -- 531	299
	 ("11111111111111111111101011110100"),	 -- 530	-1292
	 ("00000000000000000000000100101001"),	 -- 529	297
	 ("00000000000000000000000100101000"),	 -- 528	296
	 ("11111111111111111111101011111010"),	 -- 527	-1286
	 ("00000000000000000000000100100110"),	 -- 526	294
	 ("00000000000000000000000100100101"),	 -- 525	293
	 ("11111111111111111111101100000000"),	 -- 524	-1280
	 ("00000000000000000000000100100011"),	 -- 523	291
	 ("00000000000000000000000100100010"),	 -- 522	290
	 ("11111111111111111111101100000110"),	 -- 521	-1274
	 ("00000000000000000000000100100000"),	 -- 520	288
	 ("00000000000000000000000100011111"),	 -- 519	287
	 ("11111111111111111111101100001100"),	 -- 518	-1268
	 ("00000000000000000000000100011101"),	 -- 517	285
	 ("00000000000000000000000100011100"),	 -- 516	284
	 ("11111111111111111111101100010010"),	 -- 515	-1262
	 ("00000000000000000000000100011010"),	 -- 514	282
	 ("00000000000000000000000100011001"),	 -- 513	281
	 ("11111111111111111111101100011000"),	 -- 512	-1256
	 ("00000000000000000000000100010111"),	 -- 511	279
	 ("00000000000000000000000100010110"),	 -- 510	278
	 ("11111111111111111111101100011110"),	 -- 509	-1250
	 ("00000000000000000000000100010100"),	 -- 508	276
	 ("00000000000000000000000100010011"),	 -- 507	275
	 ("11111111111111111111101100100100"),	 -- 506	-1244
	 ("00000000000000000000000100010001"),	 -- 505	273
	 ("00000000000000000000000100010000"),	 -- 504	272
	 ("11111111111111111111101100101010"),	 -- 503	-1238
	 ("00000000000000000000000100001110"),	 -- 502	270
	 ("00000000000000000000000100001101"),	 -- 501	269
	 ("11111111111111111111101100110000"),	 -- 500	-1232
	 ("00000000000000000000000100001011"),	 -- 499	267
	 ("00000000000000000000000100001010"),	 -- 498	266
	 ("11111111111111111111101100110110"),	 -- 497	-1226
	 ("00000000000000000000000100001000"),	 -- 496	264
	 ("00000000000000000000000100000111"),	 -- 495	263
	 ("11111111111111111111101100111100"),	 -- 494	-1220
	 ("00000000000000000000000100000101"),	 -- 493	261
	 ("00000000000000000000000100000100"),	 -- 492	260
	 ("11111111111111111111101101000010"),	 -- 491	-1214
	 ("00000000000000000000000100000010"),	 -- 490	258
	 ("00000000000000000000000100000001"),	 -- 489	257
	 ("11111111111111111111101101001000"),	 -- 488	-1208
	 ("00000000000000000000000011111111"),	 -- 487	255
	 ("00000000000000000000000011111110"),	 -- 486	254
	 ("11111111111111111111101101001110"),	 -- 485	-1202
	 ("00000000000000000000000011111100"),	 -- 484	252
	 ("00000000000000000000000011111011"),	 -- 483	251
	 ("11111111111111111111101101010100"),	 -- 482	-1196
	 ("00000000000000000000000011111001"),	 -- 481	249
	 ("00000000000000000000000011111000"),	 -- 480	248
	 ("11111111111111111111101101011010"),	 -- 479	-1190
	 ("00000000000000000000000011110110"),	 -- 478	246
	 ("00000000000000000000000011110101"),	 -- 477	245
	 ("11111111111111111111101101100000"),	 -- 476	-1184
	 ("00000000000000000000000011110011"),	 -- 475	243
	 ("00000000000000000000000011110010"),	 -- 474	242
	 ("11111111111111111111101101100110"),	 -- 473	-1178
	 ("00000000000000000000000011110000"),	 -- 472	240
	 ("00000000000000000000000011101111"),	 -- 471	239
	 ("11111111111111111111101101101100"),	 -- 470	-1172
	 ("00000000000000000000000011101101"),	 -- 469	237
	 ("00000000000000000000000011101100"),	 -- 468	236
	 ("11111111111111111111101101110010"),	 -- 467	-1166
	 ("00000000000000000000000011101010"),	 -- 466	234
	 ("00000000000000000000000011101001"),	 -- 465	233
	 ("11111111111111111111101101111000"),	 -- 464	-1160
	 ("00000000000000000000000011100111"),	 -- 463	231
	 ("00000000000000000000000011100110"),	 -- 462	230
	 ("11111111111111111111101101111110"),	 -- 461	-1154
	 ("00000000000000000000000011100100"),	 -- 460	228
	 ("00000000000000000000000011100011"),	 -- 459	227
	 ("11111111111111111111101110000100"),	 -- 458	-1148
	 ("00000000000000000000000011100001"),	 -- 457	225
	 ("00000000000000000000000011100000"),	 -- 456	224
	 ("11111111111111111111101110001010"),	 -- 455	-1142
	 ("00000000000000000000000011011110"),	 -- 454	222
	 ("00000000000000000000000011011101"),	 -- 453	221
	 ("11111111111111111111101110010000"),	 -- 452	-1136
	 ("00000000000000000000000011011011"),	 -- 451	219
	 ("00000000000000000000000011011010"),	 -- 450	218
	 ("11111111111111111111101110010110"),	 -- 449	-1130
	 ("00000000000000000000000011011000"),	 -- 448	216
	 ("00000000000000000000000011010111"),	 -- 447	215
	 ("11111111111111111111101110011100"),	 -- 446	-1124
	 ("00000000000000000000000011010101"),	 -- 445	213
	 ("00000000000000000000000011010100"),	 -- 444	212
	 ("11111111111111111111101110100010"),	 -- 443	-1118
	 ("00000000000000000000000011010010"),	 -- 442	210
	 ("00000000000000000000000011010001"),	 -- 441	209
	 ("11111111111111111111101110101000"),	 -- 440	-1112
	 ("00000000000000000000000011001111"),	 -- 439	207
	 ("00000000000000000000000011001110"),	 -- 438	206
	 ("11111111111111111111101110101110"),	 -- 437	-1106
	 ("00000000000000000000000011001100"),	 -- 436	204
	 ("00000000000000000000000011001011"),	 -- 435	203
	 ("11111111111111111111101110110100"),	 -- 434	-1100
	 ("00000000000000000000000011001001"),	 -- 433	201
	 ("00000000000000000000000011001000"),	 -- 432	200
	 ("11111111111111111111101110111010"),	 -- 431	-1094
	 ("00000000000000000000000011000110"),	 -- 430	198
	 ("00000000000000000000000011000101"),	 -- 429	197
	 ("11111111111111111111101111000000"),	 -- 428	-1088
	 ("00000000000000000000000011000011"),	 -- 427	195
	 ("00000000000000000000000011000010"),	 -- 426	194
	 ("11111111111111111111101111000110"),	 -- 425	-1082
	 ("00000000000000000000000011000000"),	 -- 424	192
	 ("00000000000000000000000010111111"),	 -- 423	191
	 ("11111111111111111111101111001100"),	 -- 422	-1076
	 ("00000000000000000000000010111101"),	 -- 421	189
	 ("00000000000000000000000010111100"),	 -- 420	188
	 ("11111111111111111111101111010010"),	 -- 419	-1070
	 ("00000000000000000000000010111010"),	 -- 418	186
	 ("00000000000000000000000010111001"),	 -- 417	185
	 ("11111111111111111111101111011000"),	 -- 416	-1064
	 ("00000000000000000000000010110111"),	 -- 415	183
	 ("00000000000000000000000010110110"),	 -- 414	182
	 ("11111111111111111111101111011110"),	 -- 413	-1058
	 ("00000000000000000000000010110100"),	 -- 412	180
	 ("00000000000000000000000010110011"),	 -- 411	179
	 ("11111111111111111111101111100100"),	 -- 410	-1052
	 ("00000000000000000000000010110001"),	 -- 409	177
	 ("00000000000000000000000010110000"),	 -- 408	176
	 ("11111111111111111111101111101010"),	 -- 407	-1046
	 ("00000000000000000000000010101110"),	 -- 406	174
	 ("00000000000000000000000010101101"),	 -- 405	173
	 ("11111111111111111111101111110000"),	 -- 404	-1040
	 ("00000000000000000000000010101011"),	 -- 403	171
	 ("00000000000000000000000010101010"),	 -- 402	170
	 ("11111111111111111111101111110110"),	 -- 401	-1034
	 ("00000000000000000000000010101000"),	 -- 400	168
	 ("00000000000000000000000010100111"),	 -- 399	167
	 ("11111111111111111111101111111100"),	 -- 398	-1028
	 ("00000000000000000000000010100101"),	 -- 397	165
	 ("00000000000000000000000010100100"),	 -- 396	164
	 ("11111111111111111111110000000010"),	 -- 395	-1022
	 ("00000000000000000000000010100010"),	 -- 394	162
	 ("00000000000000000000000010100001"),	 -- 393	161
	 ("11111111111111111111110000001000"),	 -- 392	-1016
	 ("00000000000000000000000010011111"),	 -- 391	159
	 ("00000000000000000000000010011110"),	 -- 390	158
	 ("11111111111111111111110000001110"),	 -- 389	-1010
	 ("00000000000000000000000010011100"),	 -- 388	156
	 ("00000000000000000000000010011011"),	 -- 387	155
	 ("11111111111111111111110000010100"),	 -- 386	-1004
	 ("00000000000000000000000010011001"),	 -- 385	153
	 ("00000000000000000000000010011000"),	 -- 384	152
	 ("11111111111111111111110000011010"),	 -- 383	-998
	 ("00000000000000000000000010010110"),	 -- 382	150
	 ("00000000000000000000000010010101"),	 -- 381	149
	 ("11111111111111111111110000100000"),	 -- 380	-992
	 ("00000000000000000000000010010011"),	 -- 379	147
	 ("00000000000000000000000010010010"),	 -- 378	146
	 ("11111111111111111111110000100110"),	 -- 377	-986
	 ("00000000000000000000000010010000"),	 -- 376	144
	 ("00000000000000000000000010001111"),	 -- 375	143
	 ("11111111111111111111110000101100"),	 -- 374	-980
	 ("00000000000000000000000010001101"),	 -- 373	141
	 ("00000000000000000000000010001100"),	 -- 372	140
	 ("11111111111111111111110000110010"),	 -- 371	-974
	 ("00000000000000000000000010001010"),	 -- 370	138
	 ("00000000000000000000000010001001"),	 -- 369	137
	 ("11111111111111111111110000111000"),	 -- 368	-968
	 ("00000000000000000000000010000111"),	 -- 367	135
	 ("00000000000000000000000010000110"),	 -- 366	134
	 ("11111111111111111111110000111110"),	 -- 365	-962
	 ("00000000000000000000000010000100"),	 -- 364	132
	 ("00000000000000000000000010000011"),	 -- 363	131
	 ("11111111111111111111110001000100"),	 -- 362	-956
	 ("00000000000000000000000010000001"),	 -- 361	129
	 ("00000000000000000000000010000000"),	 -- 360	128
	 ("11111111111111111111110001001010"),	 -- 359	-950
	 ("00000000000000000000000001111110"),	 -- 358	126
	 ("00000000000000000000000001111101"),	 -- 357	125
	 ("11111111111111111111110001010000"),	 -- 356	-944
	 ("00000000000000000000000001111011"),	 -- 355	123
	 ("00000000000000000000000001111010"),	 -- 354	122
	 ("11111111111111111111110001010110"),	 -- 353	-938
	 ("00000000000000000000000001111000"),	 -- 352	120
	 ("00000000000000000000000001110111"),	 -- 351	119
	 ("11111111111111111111110001011100"),	 -- 350	-932
	 ("00000000000000000000000001110101"),	 -- 349	117
	 ("00000000000000000000000001110100"),	 -- 348	116
	 ("11111111111111111111110001100010"),	 -- 347	-926
	 ("00000000000000000000000001110010"),	 -- 346	114
	 ("00000000000000000000000001110001"),	 -- 345	113
	 ("11111111111111111111110001101000"),	 -- 344	-920
	 ("00000000000000000000000001101111"),	 -- 343	111
	 ("00000000000000000000000001101110"),	 -- 342	110
	 ("11111111111111111111110001101110"),	 -- 341	-914
	 ("00000000000000000000000001101100"),	 -- 340	108
	 ("00000000000000000000000001101011"),	 -- 339	107
	 ("11111111111111111111110001110100"),	 -- 338	-908
	 ("00000000000000000000000001101001"),	 -- 337	105
	 ("00000000000000000000000001101000"),	 -- 336	104
	 ("11111111111111111111110001111010"),	 -- 335	-902
	 ("00000000000000000000000001100110"),	 -- 334	102
	 ("00000000000000000000000001100101"),	 -- 333	101
	 ("11111111111111111111110010000000"),	 -- 332	-896
	 ("00000000000000000000000001100011"),	 -- 331	99
	 ("00000000000000000000000001100010"),	 -- 330	98
	 ("11111111111111111111110010000110"),	 -- 329	-890
	 ("00000000000000000000000001100000"),	 -- 328	96
	 ("00000000000000000000000001011111"),	 -- 327	95
	 ("11111111111111111111110010001100"),	 -- 326	-884
	 ("00000000000000000000000001011101"),	 -- 325	93
	 ("00000000000000000000000001011100"),	 -- 324	92
	 ("11111111111111111111110010010010"),	 -- 323	-878
	 ("00000000000000000000000001011010"),	 -- 322	90
	 ("00000000000000000000000001011001"),	 -- 321	89
	 ("11111111111111111111110010011000"),	 -- 320	-872
	 ("00000000000000000000000001010111"),	 -- 319	87
	 ("00000000000000000000000001010110"),	 -- 318	86
	 ("11111111111111111111110010011110"),	 -- 317	-866
	 ("00000000000000000000000001010100"),	 -- 316	84
	 ("00000000000000000000000001010011"),	 -- 315	83
	 ("11111111111111111111110010100100"),	 -- 314	-860
	 ("00000000000000000000000001010001"),	 -- 313	81
	 ("00000000000000000000000001010000"),	 -- 312	80
	 ("11111111111111111111110010101010"),	 -- 311	-854
	 ("00000000000000000000000001001110"),	 -- 310	78
	 ("00000000000000000000000001001101"),	 -- 309	77
	 ("11111111111111111111110010110000"),	 -- 308	-848
	 ("00000000000000000000000001001011"),	 -- 307	75
	 ("00000000000000000000000001001010"),	 -- 306	74
	 ("11111111111111111111110010110110"),	 -- 305	-842
	 ("00000000000000000000000001001000"),	 -- 304	72
	 ("00000000000000000000000001000111"),	 -- 303	71
	 ("11111111111111111111110010111100"),	 -- 302	-836
	 ("00000000000000000000000001000101"),	 -- 301	69
	 ("00000000000000000000000001000100"),	 -- 300	68
	 ("11111111111111111111110011000010"),	 -- 299	-830
	 ("00000000000000000000000001000010"),	 -- 298	66
	 ("00000000000000000000000001000001"),	 -- 297	65
	 ("11111111111111111111110011001000"),	 -- 296	-824
	 ("00000000000000000000000000111111"),	 -- 295	63
	 ("00000000000000000000000000111110"),	 -- 294	62
	 ("11111111111111111111110011001110"),	 -- 293	-818
	 ("00000000000000000000000000111100"),	 -- 292	60
	 ("00000000000000000000000000111011"),	 -- 291	59
	 ("11111111111111111111110011010100"),	 -- 290	-812
	 ("00000000000000000000000000111001"),	 -- 289	57
	 ("00000000000000000000000000111000"),	 -- 288	56
	 ("11111111111111111111110011011010"),	 -- 287	-806
	 ("00000000000000000000000000110110"),	 -- 286	54
	 ("00000000000000000000000000110101"),	 -- 285	53
	 ("11111111111111111111110011100000"),	 -- 284	-800
	 ("00000000000000000000000000110011"),	 -- 283	51
	 ("00000000000000000000000000110010"),	 -- 282	50
	 ("11111111111111111111110011100110"),	 -- 281	-794
	 ("00000000000000000000000000110000"),	 -- 280	48
	 ("00000000000000000000000000101111"),	 -- 279	47
	 ("11111111111111111111110011101100"),	 -- 278	-788
	 ("00000000000000000000000000101101"),	 -- 277	45
	 ("00000000000000000000000000101100"),	 -- 276	44
	 ("11111111111111111111110011110010"),	 -- 275	-782
	 ("00000000000000000000000000101010"),	 -- 274	42
	 ("00000000000000000000000000101001"),	 -- 273	41
	 ("11111111111111111111110011111000"),	 -- 272	-776
	 ("00000000000000000000000000100111"),	 -- 271	39
	 ("00000000000000000000000000100110"),	 -- 270	38
	 ("11111111111111111111110011111110"),	 -- 269	-770
	 ("00000000000000000000000000100100"),	 -- 268	36
	 ("00000000000000000000000000100011"),	 -- 267	35
	 ("11111111111111111111110100000100"),	 -- 266	-764
	 ("00000000000000000000000000100001"),	 -- 265	33
	 ("00000000000000000000000000100000"),	 -- 264	32
	 ("11111111111111111111110100001010"),	 -- 263	-758
	 ("00000000000000000000000000011110"),	 -- 262	30
	 ("00000000000000000000000000011101"),	 -- 261	29
	 ("11111111111111111111110100010000"),	 -- 260	-752
	 ("00000000000000000000000000011011"),	 -- 259	27
	 ("00000000000000000000000000011010"),	 -- 258	26
	 ("11111111111111111111110100010110"),	 -- 257	-746
	 ("00000000000000000000000000011000"),	 -- 256	24
	 ("00000000000000000000000000010111"),	 -- 255	23
	 ("11111111111111111111110100011100"),	 -- 254	-740
	 ("00000000000000000000000000010101"),	 -- 253	21
	 ("00000000000000000000000000010100"),	 -- 252	20
	 ("11111111111111111111110100100010"),	 -- 251	-734
	 ("00000000000000000000000000010010"),	 -- 250	18
	 ("00000000000000000000000000010001"),	 -- 249	17
	 ("11111111111111111111110100101000"),	 -- 248	-728
	 ("00000000000000000000000000001111"),	 -- 247	15
	 ("00000000000000000000000000001110"),	 -- 246	14
	 ("11111111111111111111110100101110"),	 -- 245	-722
	 ("00000000000000000000000000001100"),	 -- 244	12
	 ("00000000000000000000000000001011"),	 -- 243	11
	 ("11111111111111111111110100110100"),	 -- 242	-716
	 ("00000000000000000000000000001001"),	 -- 241	9
	 ("00000000000000000000000000001000"),	 -- 240	8
	 ("11111111111111111111110100111010"),	 -- 239	-710
	 ("00000000000000000000000000000110"),	 -- 238	6
	 ("00000000000000000000000000000101"),	 -- 237	5
	 ("11111111111111111111110101000000"),	 -- 236	-704
	 ("00000000000000000000000000000011"),	 -- 235	3
	 ("00000000000000000000000000000010"),	 -- 234	2
	 ("11111111111111111111110101000110"),	 -- 233	-698
	 ("00000000000000000000000000000000"),	 -- 232	0
	 ("11111111111111111111111111111111"),	 -- 231	-1
	 ("11111111111111111111110101001100"),	 -- 230	-692
	 ("11111111111111111111111111111101"),	 -- 229	-3
	 ("11111111111111111111111111111100"),	 -- 228	-4
	 ("11111111111111111111110101010010"),	 -- 227	-686
	 ("11111111111111111111111111111010"),	 -- 226	-6
	 ("11111111111111111111111111111001"),	 -- 225	-7
	 ("11111111111111111111110101011000"),	 -- 224	-680
	 ("11111111111111111111111111110111"),	 -- 223	-9
	 ("11111111111111111111111111110110"),	 -- 222	-10
	 ("11111111111111111111110101011110"),	 -- 221	-674
	 ("11111111111111111111111111110100"),	 -- 220	-12
	 ("11111111111111111111111111110011"),	 -- 219	-13
	 ("11111111111111111111110101100100"),	 -- 218	-668
	 ("11111111111111111111111111110001"),	 -- 217	-15
	 ("11111111111111111111111111110000"),	 -- 216	-16
	 ("11111111111111111111110101101010"),	 -- 215	-662
	 ("11111111111111111111111111101110"),	 -- 214	-18
	 ("11111111111111111111111111101101"),	 -- 213	-19
	 ("11111111111111111111110101110000"),	 -- 212	-656
	 ("11111111111111111111111111101011"),	 -- 211	-21
	 ("11111111111111111111111111101010"),	 -- 210	-22
	 ("11111111111111111111110101110110"),	 -- 209	-650
	 ("11111111111111111111111111101000"),	 -- 208	-24
	 ("11111111111111111111111111100111"),	 -- 207	-25
	 ("11111111111111111111110101111100"),	 -- 206	-644
	 ("11111111111111111111111111100101"),	 -- 205	-27
	 ("11111111111111111111111111100100"),	 -- 204	-28
	 ("11111111111111111111110110000010"),	 -- 203	-638
	 ("11111111111111111111111111100010"),	 -- 202	-30
	 ("11111111111111111111111111100001"),	 -- 201	-31
	 ("11111111111111111111110110001000"),	 -- 200	-632
	 ("11111111111111111111111111011111"),	 -- 199	-33
	 ("11111111111111111111111111011110"),	 -- 198	-34
	 ("11111111111111111111110110001110"),	 -- 197	-626
	 ("11111111111111111111111111011100"),	 -- 196	-36
	 ("11111111111111111111111111011011"),	 -- 195	-37
	 ("11111111111111111111110110010100"),	 -- 194	-620
	 ("11111111111111111111111111011001"),	 -- 193	-39
	 ("11111111111111111111111111011000"),	 -- 192	-40
	 ("11111111111111111111110110011010"),	 -- 191	-614
	 ("11111111111111111111111111010110"),	 -- 190	-42
	 ("11111111111111111111111111010101"),	 -- 189	-43
	 ("11111111111111111111110110100000"),	 -- 188	-608
	 ("11111111111111111111111111010011"),	 -- 187	-45
	 ("11111111111111111111111111010010"),	 -- 186	-46
	 ("11111111111111111111110110100110"),	 -- 185	-602
	 ("11111111111111111111111111010000"),	 -- 184	-48
	 ("11111111111111111111111111001111"),	 -- 183	-49
	 ("11111111111111111111110110101100"),	 -- 182	-596
	 ("11111111111111111111111111001101"),	 -- 181	-51
	 ("11111111111111111111111111001100"),	 -- 180	-52
	 ("11111111111111111111110110110010"),	 -- 179	-590
	 ("11111111111111111111111111001010"),	 -- 178	-54
	 ("11111111111111111111111111001001"),	 -- 177	-55
	 ("11111111111111111111110110111000"),	 -- 176	-584
	 ("11111111111111111111111111000111"),	 -- 175	-57
	 ("11111111111111111111111111000110"),	 -- 174	-58
	 ("11111111111111111111110110111110"),	 -- 173	-578
	 ("11111111111111111111111111000100"),	 -- 172	-60
	 ("11111111111111111111111111000011"),	 -- 171	-61
	 ("11111111111111111111110111000100"),	 -- 170	-572
	 ("11111111111111111111111111000001"),	 -- 169	-63
	 ("11111111111111111111111111000000"),	 -- 168	-64
	 ("11111111111111111111110111001010"),	 -- 167	-566
	 ("11111111111111111111111110111110"),	 -- 166	-66
	 ("11111111111111111111111110111101"),	 -- 165	-67
	 ("11111111111111111111110111010000"),	 -- 164	-560
	 ("11111111111111111111111110111011"),	 -- 163	-69
	 ("11111111111111111111111110111010"),	 -- 162	-70
	 ("11111111111111111111110111010110"),	 -- 161	-554
	 ("11111111111111111111111110111000"),	 -- 160	-72
	 ("11111111111111111111111110110111"),	 -- 159	-73
	 ("11111111111111111111110111011100"),	 -- 158	-548
	 ("11111111111111111111111110110101"),	 -- 157	-75
	 ("11111111111111111111111110110100"),	 -- 156	-76
	 ("11111111111111111111110111100010"),	 -- 155	-542
	 ("11111111111111111111111110110010"),	 -- 154	-78
	 ("11111111111111111111111110110001"),	 -- 153	-79
	 ("11111111111111111111110111101000"),	 -- 152	-536
	 ("11111111111111111111111110101111"),	 -- 151	-81
	 ("11111111111111111111111110101110"),	 -- 150	-82
	 ("11111111111111111111110111101110"),	 -- 149	-530
	 ("11111111111111111111111110101100"),	 -- 148	-84
	 ("11111111111111111111111110101011"),	 -- 147	-85
	 ("11111111111111111111110111110100"),	 -- 146	-524
	 ("11111111111111111111111110101001"),	 -- 145	-87
	 ("11111111111111111111111110101000"),	 -- 144	-88
	 ("11111111111111111111110111111010"),	 -- 143	-518
	 ("11111111111111111111111110100110"),	 -- 142	-90
	 ("11111111111111111111111110100101"),	 -- 141	-91
	 ("11111111111111111111111000000000"),	 -- 140	-512
	 ("11111111111111111111111110100011"),	 -- 139	-93
	 ("11111111111111111111111110100010"),	 -- 138	-94
	 ("11111111111111111111111000000110"),	 -- 137	-506
	 ("11111111111111111111111110100000"),	 -- 136	-96
	 ("11111111111111111111111110011111"),	 -- 135	-97
	 ("11111111111111111111111000001100"),	 -- 134	-500
	 ("11111111111111111111111110011101"),	 -- 133	-99
	 ("11111111111111111111111110011100"),	 -- 132	-100
	 ("11111111111111111111111000010010"),	 -- 131	-494
	 ("11111111111111111111111110011010"),	 -- 130	-102
	 ("11111111111111111111111110011001"),	 -- 129	-103
	 ("11111111111111111111111000011000"),	 -- 128	-488
	 ("11111111111111111111111110010111"),	 -- 127	-105
	 ("11111111111111111111111110010110"),	 -- 126	-106
	 ("11111111111111111111111000011110"),	 -- 125	-482
	 ("11111111111111111111111110010100"),	 -- 124	-108
	 ("11111111111111111111111110010011"),	 -- 123	-109
	 ("11111111111111111111111000100100"),	 -- 122	-476
	 ("11111111111111111111111110010001"),	 -- 121	-111
	 ("11111111111111111111111110010000"),	 -- 120	-112
	 ("11111111111111111111111000101010"),	 -- 119	-470
	 ("11111111111111111111111110001110"),	 -- 118	-114
	 ("11111111111111111111111110001101"),	 -- 117	-115
	 ("11111111111111111111111000110000"),	 -- 116	-464
	 ("11111111111111111111111110001011"),	 -- 115	-117
	 ("11111111111111111111111110001010"),	 -- 114	-118
	 ("11111111111111111111111000110110"),	 -- 113	-458
	 ("11111111111111111111111110001000"),	 -- 112	-120
	 ("11111111111111111111111110000111"),	 -- 111	-121
	 ("11111111111111111111111000111100"),	 -- 110	-452
	 ("11111111111111111111111110000101"),	 -- 109	-123
	 ("11111111111111111111111110000100"),	 -- 108	-124
	 ("11111111111111111111111001000010"),	 -- 107	-446
	 ("11111111111111111111111110000010"),	 -- 106	-126
	 ("11111111111111111111111110000001"),	 -- 105	-127
	 ("11111111111111111111111001001000"),	 -- 104	-440
	 ("11111111111111111111111101111111"),	 -- 103	-129
	 ("11111111111111111111111101111110"),	 -- 102	-130
	 ("11111111111111111111111001001110"),	 -- 101	-434
	 ("11111111111111111111111101111100"),	 -- 100	-132
	 ("11111111111111111111111101111011"),	 -- 99	-133
	 ("11111111111111111111111001010100"),	 -- 98	-428
	 ("11111111111111111111111101111001"),	 -- 97	-135
	 ("11111111111111111111111101111000"),	 -- 96	-136
	 ("11111111111111111111111001011010"),	 -- 95	-422
	 ("11111111111111111111111101110110"),	 -- 94	-138
	 ("11111111111111111111111101110101"),	 -- 93	-139
	 ("11111111111111111111111001100000"),	 -- 92	-416
	 ("11111111111111111111111101110011"),	 -- 91	-141
	 ("11111111111111111111111101110010"),	 -- 90	-142
	 ("11111111111111111111111001100110"),	 -- 89	-410
	 ("11111111111111111111111101110000"),	 -- 88	-144
	 ("11111111111111111111111101101111"),	 -- 87	-145
	 ("11111111111111111111111001101100"),	 -- 86	-404
	 ("11111111111111111111111101101101"),	 -- 85	-147
	 ("11111111111111111111111101101100"),	 -- 84	-148
	 ("11111111111111111111111001110010"),	 -- 83	-398
	 ("11111111111111111111111101101010"),	 -- 82	-150
	 ("11111111111111111111111101101001"),	 -- 81	-151
	 ("11111111111111111111111001111000"),	 -- 80	-392
	 ("11111111111111111111111101100111"),	 -- 79	-153
	 ("11111111111111111111111101100110"),	 -- 78	-154
	 ("11111111111111111111111001111110"),	 -- 77	-386
	 ("11111111111111111111111101100100"),	 -- 76	-156
	 ("11111111111111111111111101100011"),	 -- 75	-157
	 ("11111111111111111111111010000100"),	 -- 74	-380
	 ("11111111111111111111111101100001"),	 -- 73	-159
	 ("11111111111111111111111101100000"),	 -- 72	-160
	 ("11111111111111111111111010001010"),	 -- 71	-374
	 ("11111111111111111111111101011110"),	 -- 70	-162
	 ("11111111111111111111111101011101"),	 -- 69	-163
	 ("11111111111111111111111010010000"),	 -- 68	-368
	 ("11111111111111111111111101011011"),	 -- 67	-165
	 ("11111111111111111111111101011010"),	 -- 66	-166
	 ("11111111111111111111111010010110"),	 -- 65	-362
	 ("11111111111111111111111101011000"),	 -- 64	-168
	 ("11111111111111111111111101010111"),	 -- 63	-169
	 ("11111111111111111111111010011100"),	 -- 62	-356
	 ("11111111111111111111111101010101"),	 -- 61	-171
	 ("11111111111111111111111101010100"),	 -- 60	-172
	 ("11111111111111111111111010100010"),	 -- 59	-350
	 ("11111111111111111111111101010010"),	 -- 58	-174
	 ("11111111111111111111111101010001"),	 -- 57	-175
	 ("11111111111111111111111010101000"),	 -- 56	-344
	 ("11111111111111111111111101001111"),	 -- 55	-177
	 ("11111111111111111111111101001110"),	 -- 54	-178
	 ("11111111111111111111111010101110"),	 -- 53	-338
	 ("11111111111111111111111101001100"),	 -- 52	-180
	 ("11111111111111111111111101001011"),	 -- 51	-181
	 ("11111111111111111111111010110100"),	 -- 50	-332
	 ("11111111111111111111111101001001"),	 -- 49	-183
	 ("11111111111111111111111101001000"),	 -- 48	-184
	 ("11111111111111111111111010111010"),	 -- 47	-326
	 ("11111111111111111111111101000110"),	 -- 46	-186
	 ("11111111111111111111111101000101"),	 -- 45	-187
	 ("11111111111111111111111011000000"),	 -- 44	-320
	 ("11111111111111111111111101000011"),	 -- 43	-189
	 ("11111111111111111111111101000010"),	 -- 42	-190
	 ("11111111111111111111111011000110"),	 -- 41	-314
	 ("11111111111111111111111101000000"),	 -- 40	-192
	 ("11111111111111111111111100111111"),	 -- 39	-193
	 ("11111111111111111111111011001100"),	 -- 38	-308
	 ("11111111111111111111111100111101"),	 -- 37	-195
	 ("11111111111111111111111100111100"),	 -- 36	-196
	 ("11111111111111111111111011010010"),	 -- 35	-302
	 ("11111111111111111111111100111010"),	 -- 34	-198
	 ("11111111111111111111111100111001"),	 -- 33	-199
	 ("11111111111111111111111011011000"),	 -- 32	-296
	 ("11111111111111111111111100110111"),	 -- 31	-201
	 ("11111111111111111111111100110110"),	 -- 30	-202
	 ("11111111111111111111111011011110"),	 -- 29	-290
	 ("11111111111111111111111100110100"),	 -- 28	-204
	 ("11111111111111111111111100110011"),	 -- 27	-205
	 ("11111111111111111111111011100100"),	 -- 26	-284
	 ("11111111111111111111111100110001"),	 -- 25	-207
	 ("11111111111111111111111100110000"),	 -- 24	-208
	 ("11111111111111111111111011101010"),	 -- 23	-278
	 ("11111111111111111111111100101110"),	 -- 22	-210
	 ("11111111111111111111111100101101"),	 -- 21	-211
	 ("11111111111111111111111011110000"),	 -- 20	-272
	 ("11111111111111111111111100101011"),	 -- 19	-213
	 ("11111111111111111111111100101010"),	 -- 18	-214
	 ("11111111111111111111111011110110"),	 -- 17	-266
	 ("11111111111111111111111100101000"),	 -- 16	-216
	 ("11111111111111111111111100100111"),	 -- 15	-217
	 ("11111111111111111111111011111100"),	 -- 14	-260
	 ("11111111111111111111111100100101"),	 -- 13	-219
	 ("11111111111111111111111100100100"),	 -- 12	-220
	 ("11111111111111111111111100000010"),	 -- 11	-254
	 ("11111111111111111111111100100010"),	 -- 10	-222
	 ("11111111111111111111111100100001"),	 -- 9	-223
	 ("11111111111111111111111100001000"),	 -- 8	-248
	 ("11111111111111111111111100011111"),	 -- 7	-225
	 ("11111111111111111111111100011110"),	 -- 6	-226
	 ("11111111111111111111111100001110"),	 -- 5	-242
	 ("11111111111111111111111100011100"),	 -- 4	-228
	 ("11111111111111111111111100011011"),	 -- 3	-229
	 ("11111111111111111111111100010100"),	 -- 2	-236
	 ("11111111111111111111111100011001"),	 -- 1	-231
	 ("11111111111111111111111100011000"));	 -- 0	-232

begin
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we = '1') then
        RAM(conv_integer(address)) <= data_in;
        data_out <= RAM(conv_integer(read_a));
      elsif (oe = '1') then
        data_out <= RAM(conv_integer(read_a));
      end if;
      read_a <= address;
    end if;
  end process;
end rtl;
