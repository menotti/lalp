-- IEEE Libraries -- 
library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 

entity dual_block_ram_x is 
generic( 
	data_width : integer := 8; 
	address_width : integer := 8 
); 
port( 
	data_in_0 : in std_logic_vector(data_width-1 downto 0) := (others => '0'); 
	address_0 : in std_logic_vector(address_width-1 downto 0); 
	we_0: in std_logic := '0'; 
	oe_0: in std_logic := '1'; 
	data_out_0 : out std_logic_vector(data_width-1 downto 0); 
	data_in_1 : in std_logic_vector(data_width-1 downto 0) := (others => '0'); 
	address_1 : in std_logic_vector(address_width-1 downto 0); 
	we_1: in std_logic := '0'; 
	oe_1: in std_logic := '1'; 
	data_out_1 : out std_logic_vector(data_width-1 downto 0); 
	clk : in std_logic); 
end dual_block_ram_x; 

architecture rtl of dual_block_ram_x is 

constant mem_depth : integer := 2**address_width; 
type ram_type is array (mem_depth-1 downto 0) 
of std_logic_vector (data_width-1 downto 0); 

signal read_a : std_logic_vector(address_width-1 downto 0); 
signal read_b : std_logic_vector(address_width-1 downto 0); 
signal RAM : ram_type := ram_type'( 
	 ("00000000000000000000000000000100"),	 -- 2047	4
	 ("00000000000000000000000000000000"),	 -- 2046	0
	 ("00000000000000000000000000000000"),	 -- 2045	0
	 ("00000000000000000000000000000000"),	 -- 2044	0
	 ("00000000000000000000000000000000"),	 -- 2043	0
	 ("00000000000000000000000000000000"),	 -- 2042	0
	 ("00000000000000000000000000000000"),	 -- 2041	0
	 ("00000000000000000000000000000000"),	 -- 2040	0
	 ("00000000000000000000000000000000"),	 -- 2039	0
	 ("00000000000000000000000000000000"),	 -- 2038	0
	 ("00000000000000000000000000000000"),	 -- 2037	0
	 ("00000000000000000000000000000000"),	 -- 2036	0
	 ("00000000000000000000000000000000"),	 -- 2035	0
	 ("00000000000000000000000000000000"),	 -- 2034	0
	 ("00000000000000000000000000000000"),	 -- 2033	0
	 ("00000000000000000000000000000000"),	 -- 2032	0
	 ("00000000000000000000000000000000"),	 -- 2031	0
	 ("00000000000000000000000000000000"),	 -- 2030	0
	 ("00000000000000000000000000000000"),	 -- 2029	0
	 ("00000000000000000000000000000000"),	 -- 2028	0
	 ("00000000000000000000000000000000"),	 -- 2027	0
	 ("00000000000000000000000000000000"),	 -- 2026	0
	 ("00000000000000000000000000000000"),	 -- 2025	0
	 ("00000000000000000000000000000000"),	 -- 2024	0
	 ("00000000000000000000000000000000"),	 -- 2023	0
	 ("00000000000000000000000000000000"),	 -- 2022	0
	 ("00000000000000000000000000000000"),	 -- 2021	0
	 ("00000000000000000000000000000000"),	 -- 2020	0
	 ("00000000000000000000000000000000"),	 -- 2019	0
	 ("00000000000000000000000000000000"),	 -- 2018	0
	 ("00000000000000000000000000000000"),	 -- 2017	0
	 ("00000000000000000000000000000000"),	 -- 2016	0
	 ("00000000000000000000000000000000"),	 -- 2015	0
	 ("00000000000000000000000000000000"),	 -- 2014	0
	 ("00000000000000000000000000000000"),	 -- 2013	0
	 ("00000000000000000000000000000000"),	 -- 2012	0
	 ("00000000000000000000000000000000"),	 -- 2011	0
	 ("00000000000000000000000000000000"),	 -- 2010	0
	 ("00000000000000000000000000000000"),	 -- 2009	0
	 ("00000000000000000000000000000000"),	 -- 2008	0
	 ("00000000000000000000000000000000"),	 -- 2007	0
	 ("00000000000000000000000000000000"),	 -- 2006	0
	 ("00000000000000000000000000000000"),	 -- 2005	0
	 ("00000000000000000000000000000000"),	 -- 2004	0
	 ("00000000000000000000000000000000"),	 -- 2003	0
	 ("00000000000000000000000000000000"),	 -- 2002	0
	 ("00000000000000000000000000000000"),	 -- 2001	0
	 ("00000000000000000000000000000000"),	 -- 2000	0
	 ("00000000000000000000000000000000"),	 -- 1999	0
	 ("00000000000000000000000000000000"),	 -- 1998	0
	 ("00000000000000000000000000000000"),	 -- 1997	0
	 ("00000000000000000000000000000000"),	 -- 1996	0
	 ("00000000000000000000000000000000"),	 -- 1995	0
	 ("00000000000000000000000000000000"),	 -- 1994	0
	 ("00000000000000000000000000000000"),	 -- 1993	0
	 ("00000000000000000000000000000000"),	 -- 1992	0
	 ("00000000000000000000000000000000"),	 -- 1991	0
	 ("00000000000000000000000000000000"),	 -- 1990	0
	 ("00000000000000000000000000000000"),	 -- 1989	0
	 ("00000000000000000000000000000000"),	 -- 1988	0
	 ("00000000000000000000000000000000"),	 -- 1987	0
	 ("00000000000000000000000000000000"),	 -- 1986	0
	 ("00000000000000000000000000000000"),	 -- 1985	0
	 ("00000000000000000000000000000000"),	 -- 1984	0
	 ("00000000000000000000000000000000"),	 -- 1983	0
	 ("00000000000000000000000000000000"),	 -- 1982	0
	 ("00000000000000000000000000000000"),	 -- 1981	0
	 ("00000000000000000000000000000000"),	 -- 1980	0
	 ("00000000000000000000000000000000"),	 -- 1979	0
	 ("00000000000000000000000000000000"),	 -- 1978	0
	 ("00000000000000000000000000000000"),	 -- 1977	0
	 ("00000000000000000000000000000000"),	 -- 1976	0
	 ("00000000000000000000000000000000"),	 -- 1975	0
	 ("00000000000000000000000000000000"),	 -- 1974	0
	 ("00000000000000000000000000000000"),	 -- 1973	0
	 ("00000000000000000000000000000000"),	 -- 1972	0
	 ("00000000000000000000000000000000"),	 -- 1971	0
	 ("00000000000000000000000000000000"),	 -- 1970	0
	 ("00000000000000000000000000000000"),	 -- 1969	0
	 ("00000000000000000000000000000000"),	 -- 1968	0
	 ("00000000000000000000000000000000"),	 -- 1967	0
	 ("00000000000000000000000000000000"),	 -- 1966	0
	 ("00000000000000000000000000000000"),	 -- 1965	0
	 ("00000000000000000000000000000000"),	 -- 1964	0
	 ("00000000000000000000000000000000"),	 -- 1963	0
	 ("00000000000000000000000000000000"),	 -- 1962	0
	 ("00000000000000000000000000000000"),	 -- 1961	0
	 ("00000000000000000000000000000000"),	 -- 1960	0
	 ("00000000000000000000000000000000"),	 -- 1959	0
	 ("00000000000000000000000000000000"),	 -- 1958	0
	 ("00000000000000000000000000000000"),	 -- 1957	0
	 ("00000000000000000000000000000000"),	 -- 1956	0
	 ("00000000000000000000000000000000"),	 -- 1955	0
	 ("00000000000000000000000000000000"),	 -- 1954	0
	 ("00000000000000000000000000000000"),	 -- 1953	0
	 ("00000000000000000000000000000000"),	 -- 1952	0
	 ("00000000000000000000000000000000"),	 -- 1951	0
	 ("00000000000000000000000000000000"),	 -- 1950	0
	 ("00000000000000000000000000000000"),	 -- 1949	0
	 ("00000000000000000000000000000000"),	 -- 1948	0
	 ("00000000000000000000000000000000"),	 -- 1947	0
	 ("00000000000000000000000000000000"),	 -- 1946	0
	 ("00000000000000000000000000000000"),	 -- 1945	0
	 ("00000000000000000000000000000000"),	 -- 1944	0
	 ("00000000000000000000000000000000"),	 -- 1943	0
	 ("00000000000000000000000000000000"),	 -- 1942	0
	 ("00000000000000000000000000000000"),	 -- 1941	0
	 ("00000000000000000000000000000000"),	 -- 1940	0
	 ("00000000000000000000000000000000"),	 -- 1939	0
	 ("00000000000000000000000000000000"),	 -- 1938	0
	 ("00000000000000000000000000000000"),	 -- 1937	0
	 ("00000000000000000000000000000000"),	 -- 1936	0
	 ("00000000000000000000000000000000"),	 -- 1935	0
	 ("00000000000000000000000000000000"),	 -- 1934	0
	 ("00000000000000000000000000000000"),	 -- 1933	0
	 ("00000000000000000000000000000000"),	 -- 1932	0
	 ("00000000000000000000000000000000"),	 -- 1931	0
	 ("00000000000000000000000000000000"),	 -- 1930	0
	 ("00000000000000000000000000000000"),	 -- 1929	0
	 ("00000000000000000000000000000000"),	 -- 1928	0
	 ("00000000000000000000000000000000"),	 -- 1927	0
	 ("00000000000000000000000000000000"),	 -- 1926	0
	 ("00000000000000000000000000000000"),	 -- 1925	0
	 ("00000000000000000000000000000000"),	 -- 1924	0
	 ("00000000000000000000000000000000"),	 -- 1923	0
	 ("00000000000000000000000000000000"),	 -- 1922	0
	 ("00000000000000000000000000000000"),	 -- 1921	0
	 ("00000000000000000000000000000000"),	 -- 1920	0
	 ("00000000000000000000000000000000"),	 -- 1919	0
	 ("00000000000000000000000000000000"),	 -- 1918	0
	 ("00000000000000000000000000000000"),	 -- 1917	0
	 ("00000000000000000000000000000000"),	 -- 1916	0
	 ("00000000000000000000000000000000"),	 -- 1915	0
	 ("00000000000000000000000000000000"),	 -- 1914	0
	 ("00000000000000000000000000000000"),	 -- 1913	0
	 ("00000000000000000000000000000000"),	 -- 1912	0
	 ("00000000000000000000000000000000"),	 -- 1911	0
	 ("00000000000000000000000000000000"),	 -- 1910	0
	 ("00000000000000000000000000000000"),	 -- 1909	0
	 ("00000000000000000000000000000000"),	 -- 1908	0
	 ("00000000000000000000000000000000"),	 -- 1907	0
	 ("00000000000000000000000000000000"),	 -- 1906	0
	 ("00000000000000000000000000000000"),	 -- 1905	0
	 ("00000000000000000000000000000000"),	 -- 1904	0
	 ("00000000000000000000000000000000"),	 -- 1903	0
	 ("00000000000000000000000000000000"),	 -- 1902	0
	 ("00000000000000000000000000000000"),	 -- 1901	0
	 ("00000000000000000000000000000000"),	 -- 1900	0
	 ("00000000000000000000000000000000"),	 -- 1899	0
	 ("00000000000000000000000000000000"),	 -- 1898	0
	 ("00000000000000000000000000000000"),	 -- 1897	0
	 ("00000000000000000000000000000000"),	 -- 1896	0
	 ("00000000000000000000000000000000"),	 -- 1895	0
	 ("00000000000000000000000000000000"),	 -- 1894	0
	 ("00000000000000000000000000000000"),	 -- 1893	0
	 ("00000000000000000000000000000000"),	 -- 1892	0
	 ("00000000000000000000000000000000"),	 -- 1891	0
	 ("00000000000000000000000000000000"),	 -- 1890	0
	 ("00000000000000000000000000000000"),	 -- 1889	0
	 ("00000000000000000000000000000000"),	 -- 1888	0
	 ("00000000000000000000000000000000"),	 -- 1887	0
	 ("00000000000000000000000000000000"),	 -- 1886	0
	 ("00000000000000000000000000000000"),	 -- 1885	0
	 ("00000000000000000000000000000000"),	 -- 1884	0
	 ("00000000000000000000000000000000"),	 -- 1883	0
	 ("00000000000000000000000000000000"),	 -- 1882	0
	 ("00000000000000000000000000000000"),	 -- 1881	0
	 ("00000000000000000000000000000000"),	 -- 1880	0
	 ("00000000000000000000000000000000"),	 -- 1879	0
	 ("00000000000000000000000000000000"),	 -- 1878	0
	 ("00000000000000000000000000000000"),	 -- 1877	0
	 ("00000000000000000000000000000000"),	 -- 1876	0
	 ("00000000000000000000000000000000"),	 -- 1875	0
	 ("00000000000000000000000000000000"),	 -- 1874	0
	 ("00000000000000000000000000000000"),	 -- 1873	0
	 ("00000000000000000000000000000000"),	 -- 1872	0
	 ("00000000000000000000000000000000"),	 -- 1871	0
	 ("00000000000000000000000000000000"),	 -- 1870	0
	 ("00000000000000000000000000000000"),	 -- 1869	0
	 ("00000000000000000000000000000000"),	 -- 1868	0
	 ("00000000000000000000000000000000"),	 -- 1867	0
	 ("00000000000000000000000000000000"),	 -- 1866	0
	 ("00000000000000000000000000000000"),	 -- 1865	0
	 ("00000000000000000000000000000000"),	 -- 1864	0
	 ("00000000000000000000000000000000"),	 -- 1863	0
	 ("00000000000000000000000000000000"),	 -- 1862	0
	 ("00000000000000000000000000000000"),	 -- 1861	0
	 ("00000000000000000000000000000000"),	 -- 1860	0
	 ("00000000000000000000000000000000"),	 -- 1859	0
	 ("00000000000000000000000000000000"),	 -- 1858	0
	 ("00000000000000000000000000000000"),	 -- 1857	0
	 ("00000000000000000000000000000000"),	 -- 1856	0
	 ("00000000000000000000000000000000"),	 -- 1855	0
	 ("00000000000000000000000000000000"),	 -- 1854	0
	 ("00000000000000000000000000000000"),	 -- 1853	0
	 ("00000000000000000000000000000000"),	 -- 1852	0
	 ("00000000000000000000000000000000"),	 -- 1851	0
	 ("00000000000000000000000000000000"),	 -- 1850	0
	 ("00000000000000000000000000000000"),	 -- 1849	0
	 ("00000000000000000000000000000000"),	 -- 1848	0
	 ("00000000000000000000000000000000"),	 -- 1847	0
	 ("00000000000000000000000000000000"),	 -- 1846	0
	 ("00000000000000000000000000000000"),	 -- 1845	0
	 ("00000000000000000000000000000000"),	 -- 1844	0
	 ("00000000000000000000000000000000"),	 -- 1843	0
	 ("00000000000000000000000000000000"),	 -- 1842	0
	 ("00000000000000000000000000000000"),	 -- 1841	0
	 ("00000000000000000000000000000000"),	 -- 1840	0
	 ("00000000000000000000000000000000"),	 -- 1839	0
	 ("00000000000000000000000000000000"),	 -- 1838	0
	 ("00000000000000000000000000000000"),	 -- 1837	0
	 ("00000000000000000000000000000000"),	 -- 1836	0
	 ("00000000000000000000000000000000"),	 -- 1835	0
	 ("00000000000000000000000000000000"),	 -- 1834	0
	 ("00000000000000000000000000000000"),	 -- 1833	0
	 ("00000000000000000000000000000000"),	 -- 1832	0
	 ("00000000000000000000000000000000"),	 -- 1831	0
	 ("00000000000000000000000000000000"),	 -- 1830	0
	 ("00000000000000000000000000000000"),	 -- 1829	0
	 ("00000000000000000000000000000000"),	 -- 1828	0
	 ("00000000000000000000000000000000"),	 -- 1827	0
	 ("00000000000000000000000000000000"),	 -- 1826	0
	 ("00000000000000000000000000000000"),	 -- 1825	0
	 ("00000000000000000000000000000000"),	 -- 1824	0
	 ("00000000000000000000000000000000"),	 -- 1823	0
	 ("00000000000000000000000000000000"),	 -- 1822	0
	 ("00000000000000000000000000000000"),	 -- 1821	0
	 ("00000000000000000000000000000000"),	 -- 1820	0
	 ("00000000000000000000000000000000"),	 -- 1819	0
	 ("00000000000000000000000000000000"),	 -- 1818	0
	 ("00000000000000000000000000000000"),	 -- 1817	0
	 ("00000000000000000000000000000000"),	 -- 1816	0
	 ("00000000000000000000000000000000"),	 -- 1815	0
	 ("00000000000000000000000000000000"),	 -- 1814	0
	 ("00000000000000000000000000000000"),	 -- 1813	0
	 ("00000000000000000000000000000000"),	 -- 1812	0
	 ("00000000000000000000000000000000"),	 -- 1811	0
	 ("00000000000000000000000000000000"),	 -- 1810	0
	 ("00000000000000000000000000000000"),	 -- 1809	0
	 ("00000000000000000000000000000000"),	 -- 1808	0
	 ("00000000000000000000000000000000"),	 -- 1807	0
	 ("00000000000000000000000000000000"),	 -- 1806	0
	 ("00000000000000000000000000000000"),	 -- 1805	0
	 ("00000000000000000000000000000000"),	 -- 1804	0
	 ("00000000000000000000000000000000"),	 -- 1803	0
	 ("00000000000000000000000000000000"),	 -- 1802	0
	 ("00000000000000000000000000000000"),	 -- 1801	0
	 ("00000000000000000000000000000000"),	 -- 1800	0
	 ("00000000000000000000000000000000"),	 -- 1799	0
	 ("00000000000000000000000000000000"),	 -- 1798	0
	 ("00000000000000000000000000000000"),	 -- 1797	0
	 ("00000000000000000000000000000000"),	 -- 1796	0
	 ("00000000000000000000000000000000"),	 -- 1795	0
	 ("00000000000000000000000000000000"),	 -- 1794	0
	 ("00000000000000000000000000000000"),	 -- 1793	0
	 ("00000000000000000000000000000000"),	 -- 1792	0
	 ("00000000000000000000000000000000"),	 -- 1791	0
	 ("00000000000000000000000000000000"),	 -- 1790	0
	 ("00000000000000000000000000000000"),	 -- 1789	0
	 ("00000000000000000000000000000000"),	 -- 1788	0
	 ("00000000000000000000000000000000"),	 -- 1787	0
	 ("00000000000000000000000000000000"),	 -- 1786	0
	 ("00000000000000000000000000000000"),	 -- 1785	0
	 ("00000000000000000000000000000000"),	 -- 1784	0
	 ("00000000000000000000000000000000"),	 -- 1783	0
	 ("00000000000000000000000000000000"),	 -- 1782	0
	 ("00000000000000000000000000000000"),	 -- 1781	0
	 ("00000000000000000000000000000000"),	 -- 1780	0
	 ("00000000000000000000000000000000"),	 -- 1779	0
	 ("00000000000000000000000000000000"),	 -- 1778	0
	 ("00000000000000000000000000000000"),	 -- 1777	0
	 ("00000000000000000000000000000000"),	 -- 1776	0
	 ("00000000000000000000000000000000"),	 -- 1775	0
	 ("00000000000000000000000000000000"),	 -- 1774	0
	 ("00000000000000000000000000000000"),	 -- 1773	0
	 ("00000000000000000000000000000000"),	 -- 1772	0
	 ("00000000000000000000000000000000"),	 -- 1771	0
	 ("00000000000000000000000000000000"),	 -- 1770	0
	 ("00000000000000000000000000000000"),	 -- 1769	0
	 ("00000000000000000000000000000000"),	 -- 1768	0
	 ("00000000000000000000000000000000"),	 -- 1767	0
	 ("00000000000000000000000000000000"),	 -- 1766	0
	 ("00000000000000000000000000000000"),	 -- 1765	0
	 ("00000000000000000000000000000000"),	 -- 1764	0
	 ("00000000000000000000000000000000"),	 -- 1763	0
	 ("00000000000000000000000000000000"),	 -- 1762	0
	 ("00000000000000000000000000000000"),	 -- 1761	0
	 ("00000000000000000000000000000000"),	 -- 1760	0
	 ("00000000000000000000000000000000"),	 -- 1759	0
	 ("00000000000000000000000000000000"),	 -- 1758	0
	 ("00000000000000000000000000000000"),	 -- 1757	0
	 ("00000000000000000000000000000000"),	 -- 1756	0
	 ("00000000000000000000000000000000"),	 -- 1755	0
	 ("00000000000000000000000000000000"),	 -- 1754	0
	 ("00000000000000000000000000000000"),	 -- 1753	0
	 ("00000000000000000000000000000000"),	 -- 1752	0
	 ("00000000000000000000000000000000"),	 -- 1751	0
	 ("00000000000000000000000000000000"),	 -- 1750	0
	 ("00000000000000000000000000000000"),	 -- 1749	0
	 ("00000000000000000000000000000000"),	 -- 1748	0
	 ("00000000000000000000000000000000"),	 -- 1747	0
	 ("00000000000000000000000000000000"),	 -- 1746	0
	 ("00000000000000000000000000000000"),	 -- 1745	0
	 ("00000000000000000000000000000000"),	 -- 1744	0
	 ("00000000000000000000000000000000"),	 -- 1743	0
	 ("00000000000000000000000000000000"),	 -- 1742	0
	 ("00000000000000000000000000000000"),	 -- 1741	0
	 ("00000000000000000000000000000000"),	 -- 1740	0
	 ("00000000000000000000000000000000"),	 -- 1739	0
	 ("00000000000000000000000000000000"),	 -- 1738	0
	 ("00000000000000000000000000000000"),	 -- 1737	0
	 ("00000000000000000000000000000000"),	 -- 1736	0
	 ("00000000000000000000000000000000"),	 -- 1735	0
	 ("00000000000000000000000000000000"),	 -- 1734	0
	 ("00000000000000000000000000000000"),	 -- 1733	0
	 ("00000000000000000000000000000000"),	 -- 1732	0
	 ("00000000000000000000000000000000"),	 -- 1731	0
	 ("00000000000000000000000000000000"),	 -- 1730	0
	 ("00000000000000000000000000000000"),	 -- 1729	0
	 ("00000000000000000000000000000000"),	 -- 1728	0
	 ("00000000000000000000000000000000"),	 -- 1727	0
	 ("00000000000000000000000000000000"),	 -- 1726	0
	 ("00000000000000000000000000000000"),	 -- 1725	0
	 ("00000000000000000000000000000000"),	 -- 1724	0
	 ("00000000000000000000000000000000"),	 -- 1723	0
	 ("00000000000000000000000000000000"),	 -- 1722	0
	 ("00000000000000000000000000000000"),	 -- 1721	0
	 ("00000000000000000000000000000000"),	 -- 1720	0
	 ("00000000000000000000000000000000"),	 -- 1719	0
	 ("00000000000000000000000000000000"),	 -- 1718	0
	 ("00000000000000000000000000000000"),	 -- 1717	0
	 ("00000000000000000000000000000000"),	 -- 1716	0
	 ("00000000000000000000000000000000"),	 -- 1715	0
	 ("00000000000000000000000000000000"),	 -- 1714	0
	 ("00000000000000000000000000000000"),	 -- 1713	0
	 ("00000000000000000000000000000000"),	 -- 1712	0
	 ("00000000000000000000000000000000"),	 -- 1711	0
	 ("00000000000000000000000000000000"),	 -- 1710	0
	 ("00000000000000000000000000000000"),	 -- 1709	0
	 ("00000000000000000000000000000000"),	 -- 1708	0
	 ("00000000000000000000000000000000"),	 -- 1707	0
	 ("00000000000000000000000000000000"),	 -- 1706	0
	 ("00000000000000000000000000000000"),	 -- 1705	0
	 ("00000000000000000000000000000000"),	 -- 1704	0
	 ("00000000000000000000000000000000"),	 -- 1703	0
	 ("00000000000000000000000000000000"),	 -- 1702	0
	 ("00000000000000000000000000000000"),	 -- 1701	0
	 ("00000000000000000000000000000000"),	 -- 1700	0
	 ("00000000000000000000000000000000"),	 -- 1699	0
	 ("00000000000000000000000000000000"),	 -- 1698	0
	 ("00000000000000000000000000000000"),	 -- 1697	0
	 ("00000000000000000000000000000000"),	 -- 1696	0
	 ("00000000000000000000000000000000"),	 -- 1695	0
	 ("00000000000000000000000000000000"),	 -- 1694	0
	 ("00000000000000000000000000000000"),	 -- 1693	0
	 ("00000000000000000000000000000000"),	 -- 1692	0
	 ("00000000000000000000000000000000"),	 -- 1691	0
	 ("00000000000000000000000000000000"),	 -- 1690	0
	 ("00000000000000000000000000000000"),	 -- 1689	0
	 ("00000000000000000000000000000000"),	 -- 1688	0
	 ("00000000000000000000000000000000"),	 -- 1687	0
	 ("00000000000000000000000000000000"),	 -- 1686	0
	 ("00000000000000000000000000000000"),	 -- 1685	0
	 ("00000000000000000000000000000000"),	 -- 1684	0
	 ("00000000000000000000000000000000"),	 -- 1683	0
	 ("00000000000000000000000000000000"),	 -- 1682	0
	 ("00000000000000000000000000000000"),	 -- 1681	0
	 ("00000000000000000000000000000000"),	 -- 1680	0
	 ("00000000000000000000000000000000"),	 -- 1679	0
	 ("00000000000000000000000000000000"),	 -- 1678	0
	 ("00000000000000000000000000000000"),	 -- 1677	0
	 ("00000000000000000000000000000000"),	 -- 1676	0
	 ("00000000000000000000000000000000"),	 -- 1675	0
	 ("00000000000000000000000000000000"),	 -- 1674	0
	 ("00000000000000000000000000000000"),	 -- 1673	0
	 ("00000000000000000000000000000000"),	 -- 1672	0
	 ("00000000000000000000000000000000"),	 -- 1671	0
	 ("00000000000000000000000000000000"),	 -- 1670	0
	 ("00000000000000000000000000000000"),	 -- 1669	0
	 ("00000000000000000000000000000000"),	 -- 1668	0
	 ("00000000000000000000000000000000"),	 -- 1667	0
	 ("00000000000000000000000000000000"),	 -- 1666	0
	 ("00000000000000000000000000000000"),	 -- 1665	0
	 ("00000000000000000000000000000000"),	 -- 1664	0
	 ("00000000000000000000000000000000"),	 -- 1663	0
	 ("00000000000000000000000000000000"),	 -- 1662	0
	 ("00000000000000000000000000000000"),	 -- 1661	0
	 ("00000000000000000000000000000000"),	 -- 1660	0
	 ("00000000000000000000000000000000"),	 -- 1659	0
	 ("00000000000000000000000000000000"),	 -- 1658	0
	 ("00000000000000000000000000000000"),	 -- 1657	0
	 ("00000000000000000000000000000000"),	 -- 1656	0
	 ("00000000000000000000000000000000"),	 -- 1655	0
	 ("00000000000000000000000000000000"),	 -- 1654	0
	 ("00000000000000000000000000000000"),	 -- 1653	0
	 ("00000000000000000000000000000000"),	 -- 1652	0
	 ("00000000000000000000000000000000"),	 -- 1651	0
	 ("00000000000000000000000000000000"),	 -- 1650	0
	 ("00000000000000000000000000000000"),	 -- 1649	0
	 ("00000000000000000000000000000000"),	 -- 1648	0
	 ("00000000000000000000000000000000"),	 -- 1647	0
	 ("00000000000000000000000000000000"),	 -- 1646	0
	 ("00000000000000000000000000000000"),	 -- 1645	0
	 ("00000000000000000000000000000000"),	 -- 1644	0
	 ("00000000000000000000000000000000"),	 -- 1643	0
	 ("00000000000000000000000000000000"),	 -- 1642	0
	 ("00000000000000000000000000000000"),	 -- 1641	0
	 ("00000000000000000000000000000000"),	 -- 1640	0
	 ("00000000000000000000000000000000"),	 -- 1639	0
	 ("00000000000000000000000000000000"),	 -- 1638	0
	 ("00000000000000000000000000000000"),	 -- 1637	0
	 ("00000000000000000000000000000000"),	 -- 1636	0
	 ("00000000000000000000000000000000"),	 -- 1635	0
	 ("00000000000000000000000000000000"),	 -- 1634	0
	 ("00000000000000000000000000000000"),	 -- 1633	0
	 ("00000000000000000000000000000000"),	 -- 1632	0
	 ("00000000000000000000000000000000"),	 -- 1631	0
	 ("00000000000000000000000000000000"),	 -- 1630	0
	 ("00000000000000000000000000000000"),	 -- 1629	0
	 ("00000000000000000000000000000000"),	 -- 1628	0
	 ("00000000000000000000000000000000"),	 -- 1627	0
	 ("00000000000000000000000000000000"),	 -- 1626	0
	 ("00000000000000000000000000000000"),	 -- 1625	0
	 ("00000000000000000000000000000000"),	 -- 1624	0
	 ("00000000000000000000000000000000"),	 -- 1623	0
	 ("00000000000000000000000000000000"),	 -- 1622	0
	 ("00000000000000000000000000000000"),	 -- 1621	0
	 ("00000000000000000000000000000000"),	 -- 1620	0
	 ("00000000000000000000000000000000"),	 -- 1619	0
	 ("00000000000000000000000000000000"),	 -- 1618	0
	 ("00000000000000000000000000000000"),	 -- 1617	0
	 ("00000000000000000000000000000000"),	 -- 1616	0
	 ("00000000000000000000000000000000"),	 -- 1615	0
	 ("00000000000000000000000000000000"),	 -- 1614	0
	 ("00000000000000000000000000000000"),	 -- 1613	0
	 ("00000000000000000000000000000000"),	 -- 1612	0
	 ("00000000000000000000000000000000"),	 -- 1611	0
	 ("00000000000000000000000000000000"),	 -- 1610	0
	 ("00000000000000000000000000000000"),	 -- 1609	0
	 ("00000000000000000000000000000000"),	 -- 1608	0
	 ("00000000000000000000000000000000"),	 -- 1607	0
	 ("00000000000000000000000000000000"),	 -- 1606	0
	 ("00000000000000000000000000000000"),	 -- 1605	0
	 ("00000000000000000000000000000000"),	 -- 1604	0
	 ("00000000000000000000000000000000"),	 -- 1603	0
	 ("00000000000000000000000000000000"),	 -- 1602	0
	 ("00000000000000000000000000000000"),	 -- 1601	0
	 ("00000000000000000000000000000000"),	 -- 1600	0
	 ("00000000000000000000000000000000"),	 -- 1599	0
	 ("00000000000000000000000000000000"),	 -- 1598	0
	 ("00000000000000000000000000000000"),	 -- 1597	0
	 ("00000000000000000000000000000000"),	 -- 1596	0
	 ("00000000000000000000000000000000"),	 -- 1595	0
	 ("00000000000000000000000000000000"),	 -- 1594	0
	 ("00000000000000000000000000000000"),	 -- 1593	0
	 ("00000000000000000000000000000000"),	 -- 1592	0
	 ("00000000000000000000000000000000"),	 -- 1591	0
	 ("00000000000000000000000000000000"),	 -- 1590	0
	 ("00000000000000000000000000000000"),	 -- 1589	0
	 ("00000000000000000000000000000000"),	 -- 1588	0
	 ("00000000000000000000000000000000"),	 -- 1587	0
	 ("00000000000000000000000000000000"),	 -- 1586	0
	 ("00000000000000000000000000000000"),	 -- 1585	0
	 ("00000000000000000000000000000000"),	 -- 1584	0
	 ("00000000000000000000000000000000"),	 -- 1583	0
	 ("00000000000000000000000000000000"),	 -- 1582	0
	 ("00000000000000000000000000000000"),	 -- 1581	0
	 ("00000000000000000000000000000000"),	 -- 1580	0
	 ("00000000000000000000000000000000"),	 -- 1579	0
	 ("00000000000000000000000000000000"),	 -- 1578	0
	 ("00000000000000000000000000000000"),	 -- 1577	0
	 ("00000000000000000000000000000000"),	 -- 1576	0
	 ("00000000000000000000000000000000"),	 -- 1575	0
	 ("00000000000000000000000000000000"),	 -- 1574	0
	 ("00000000000000000000000000000000"),	 -- 1573	0
	 ("00000000000000000000000000000000"),	 -- 1572	0
	 ("00000000000000000000000000000000"),	 -- 1571	0
	 ("00000000000000000000000000000000"),	 -- 1570	0
	 ("00000000000000000000000000000000"),	 -- 1569	0
	 ("00000000000000000000000000000000"),	 -- 1568	0
	 ("00000000000000000000000000000000"),	 -- 1567	0
	 ("00000000000000000000000000000000"),	 -- 1566	0
	 ("00000000000000000000000000000000"),	 -- 1565	0
	 ("00000000000000000000000000000000"),	 -- 1564	0
	 ("00000000000000000000000000000000"),	 -- 1563	0
	 ("00000000000000000000000000000000"),	 -- 1562	0
	 ("00000000000000000000000000000000"),	 -- 1561	0
	 ("00000000000000000000000000000000"),	 -- 1560	0
	 ("00000000000000000000000000000000"),	 -- 1559	0
	 ("00000000000000000000000000000000"),	 -- 1558	0
	 ("00000000000000000000000000000000"),	 -- 1557	0
	 ("00000000000000000000000000000000"),	 -- 1556	0
	 ("00000000000000000000000000000000"),	 -- 1555	0
	 ("00000000000000000000000000000000"),	 -- 1554	0
	 ("00000000000000000000000000000000"),	 -- 1553	0
	 ("00000000000000000000000000000000"),	 -- 1552	0
	 ("00000000000000000000000000000000"),	 -- 1551	0
	 ("00000000000000000000000000000000"),	 -- 1550	0
	 ("00000000000000000000000000000000"),	 -- 1549	0
	 ("00000000000000000000000000000000"),	 -- 1548	0
	 ("00000000000000000000000000000000"),	 -- 1547	0
	 ("00000000000000000000000000000000"),	 -- 1546	0
	 ("00000000000000000000000000000000"),	 -- 1545	0
	 ("00000000000000000000000000000000"),	 -- 1544	0
	 ("00000000000000000000000000000000"),	 -- 1543	0
	 ("00000000000000000000000000000000"),	 -- 1542	0
	 ("00000000000000000000000000000000"),	 -- 1541	0
	 ("00000000000000000000000000000000"),	 -- 1540	0
	 ("00000000000000000000000000000000"),	 -- 1539	0
	 ("00000000000000000000000000000000"),	 -- 1538	0
	 ("00000000000000000000000000000000"),	 -- 1537	0
	 ("00000000000000000000000000000000"),	 -- 1536	0
	 ("00000000000000000000000000000000"),	 -- 1535	0
	 ("00000000000000000000000000000000"),	 -- 1534	0
	 ("00000000000000000000000000000000"),	 -- 1533	0
	 ("00000000000000000000000000000000"),	 -- 1532	0
	 ("00000000000000000000000000000000"),	 -- 1531	0
	 ("00000000000000000000000000000000"),	 -- 1530	0
	 ("00000000000000000000000000000000"),	 -- 1529	0
	 ("00000000000000000000000000000000"),	 -- 1528	0
	 ("00000000000000000000000000000000"),	 -- 1527	0
	 ("00000000000000000000000000000000"),	 -- 1526	0
	 ("00000000000000000000000000000000"),	 -- 1525	0
	 ("00000000000000000000000000000000"),	 -- 1524	0
	 ("00000000000000000000000000000000"),	 -- 1523	0
	 ("00000000000000000000000000000000"),	 -- 1522	0
	 ("00000000000000000000000000000000"),	 -- 1521	0
	 ("00000000000000000000000000000000"),	 -- 1520	0
	 ("00000000000000000000000000000000"),	 -- 1519	0
	 ("00000000000000000000000000000000"),	 -- 1518	0
	 ("00000000000000000000000000000000"),	 -- 1517	0
	 ("00000000000000000000000000000000"),	 -- 1516	0
	 ("00000000000000000000000000000000"),	 -- 1515	0
	 ("00000000000000000000000000000000"),	 -- 1514	0
	 ("00000000000000000000000000000000"),	 -- 1513	0
	 ("00000000000000000000000000000000"),	 -- 1512	0
	 ("00000000000000000000000000000000"),	 -- 1511	0
	 ("00000000000000000000000000000000"),	 -- 1510	0
	 ("00000000000000000000000000000000"),	 -- 1509	0
	 ("00000000000000000000000000000000"),	 -- 1508	0
	 ("00000000000000000000000000000000"),	 -- 1507	0
	 ("00000000000000000000000000000000"),	 -- 1506	0
	 ("00000000000000000000000000000000"),	 -- 1505	0
	 ("00000000000000000000000000000000"),	 -- 1504	0
	 ("00000000000000000000000000000000"),	 -- 1503	0
	 ("00000000000000000000000000000000"),	 -- 1502	0
	 ("00000000000000000000000000000000"),	 -- 1501	0
	 ("00000000000000000000000000000000"),	 -- 1500	0
	 ("00000000000000000000000000000000"),	 -- 1499	0
	 ("00000000000000000000000000000000"),	 -- 1498	0
	 ("00000000000000000000000000000000"),	 -- 1497	0
	 ("00000000000000000000000000000000"),	 -- 1496	0
	 ("00000000000000000000000000000000"),	 -- 1495	0
	 ("00000000000000000000000000000000"),	 -- 1494	0
	 ("00000000000000000000000000000000"),	 -- 1493	0
	 ("00000000000000000000000000000000"),	 -- 1492	0
	 ("00000000000000000000000000000000"),	 -- 1491	0
	 ("00000000000000000000000000000000"),	 -- 1490	0
	 ("00000000000000000000000000000000"),	 -- 1489	0
	 ("00000000000000000000000000000000"),	 -- 1488	0
	 ("00000000000000000000000000000000"),	 -- 1487	0
	 ("00000000000000000000000000000000"),	 -- 1486	0
	 ("00000000000000000000000000000000"),	 -- 1485	0
	 ("00000000000000000000000000000000"),	 -- 1484	0
	 ("00000000000000000000000000000000"),	 -- 1483	0
	 ("00000000000000000000000000000000"),	 -- 1482	0
	 ("00000000000000000000000000000000"),	 -- 1481	0
	 ("00000000000000000000000000000000"),	 -- 1480	0
	 ("00000000000000000000000000000000"),	 -- 1479	0
	 ("00000000000000000000000000000000"),	 -- 1478	0
	 ("00000000000000000000000000000000"),	 -- 1477	0
	 ("00000000000000000000000000000000"),	 -- 1476	0
	 ("00000000000000000000000000000000"),	 -- 1475	0
	 ("00000000000000000000000000000000"),	 -- 1474	0
	 ("00000000000000000000000000000000"),	 -- 1473	0
	 ("00000000000000000000000000000000"),	 -- 1472	0
	 ("00000000000000000000000000000000"),	 -- 1471	0
	 ("00000000000000000000000000000000"),	 -- 1470	0
	 ("00000000000000000000000000000000"),	 -- 1469	0
	 ("00000000000000000000000000000000"),	 -- 1468	0
	 ("00000000000000000000000000000000"),	 -- 1467	0
	 ("00000000000000000000000000000000"),	 -- 1466	0
	 ("00000000000000000000000000000000"),	 -- 1465	0
	 ("00000000000000000000000000000000"),	 -- 1464	0
	 ("00000000000000000000000000000000"),	 -- 1463	0
	 ("00000000000000000000000000000000"),	 -- 1462	0
	 ("00000000000000000000000000000000"),	 -- 1461	0
	 ("00000000000000000000000000000000"),	 -- 1460	0
	 ("00000000000000000000000000000000"),	 -- 1459	0
	 ("00000000000000000000000000000000"),	 -- 1458	0
	 ("00000000000000000000000000000000"),	 -- 1457	0
	 ("00000000000000000000000000000000"),	 -- 1456	0
	 ("00000000000000000000000000000000"),	 -- 1455	0
	 ("00000000000000000000000000000000"),	 -- 1454	0
	 ("00000000000000000000000000000000"),	 -- 1453	0
	 ("00000000000000000000000000000000"),	 -- 1452	0
	 ("00000000000000000000000000000000"),	 -- 1451	0
	 ("00000000000000000000000000000000"),	 -- 1450	0
	 ("00000000000000000000000000000000"),	 -- 1449	0
	 ("00000000000000000000000000000000"),	 -- 1448	0
	 ("00000000000000000000000000000000"),	 -- 1447	0
	 ("00000000000000000000000000000000"),	 -- 1446	0
	 ("00000000000000000000000000000000"),	 -- 1445	0
	 ("00000000000000000000000000000000"),	 -- 1444	0
	 ("00000000000000000000000000000000"),	 -- 1443	0
	 ("00000000000000000000000000000000"),	 -- 1442	0
	 ("00000000000000000000000000000000"),	 -- 1441	0
	 ("00000000000000000000000000000000"),	 -- 1440	0
	 ("00000000000000000000000000000000"),	 -- 1439	0
	 ("00000000000000000000000000000000"),	 -- 1438	0
	 ("00000000000000000000000000000000"),	 -- 1437	0
	 ("00000000000000000000000000000000"),	 -- 1436	0
	 ("00000000000000000000000000000000"),	 -- 1435	0
	 ("00000000000000000000000000000000"),	 -- 1434	0
	 ("00000000000000000000000000000000"),	 -- 1433	0
	 ("00000000000000000000000000000000"),	 -- 1432	0
	 ("00000000000000000000000000000000"),	 -- 1431	0
	 ("00000000000000000000000000000000"),	 -- 1430	0
	 ("00000000000000000000000000000000"),	 -- 1429	0
	 ("00000000000000000000000000000000"),	 -- 1428	0
	 ("00000000000000000000000000000000"),	 -- 1427	0
	 ("00000000000000000000000000000000"),	 -- 1426	0
	 ("00000000000000000000000000000000"),	 -- 1425	0
	 ("00000000000000000000000000000000"),	 -- 1424	0
	 ("00000000000000000000000000000000"),	 -- 1423	0
	 ("00000000000000000000000000000000"),	 -- 1422	0
	 ("00000000000000000000000000000000"),	 -- 1421	0
	 ("00000000000000000000000000000000"),	 -- 1420	0
	 ("00000000000000000000000000000000"),	 -- 1419	0
	 ("00000000000000000000000000000000"),	 -- 1418	0
	 ("00000000000000000000000000000000"),	 -- 1417	0
	 ("00000000000000000000000000000000"),	 -- 1416	0
	 ("00000000000000000000000000000000"),	 -- 1415	0
	 ("00000000000000000000000000000000"),	 -- 1414	0
	 ("00000000000000000000000000000000"),	 -- 1413	0
	 ("00000000000000000000000000000000"),	 -- 1412	0
	 ("00000000000000000000000000000000"),	 -- 1411	0
	 ("00000000000000000000000000000000"),	 -- 1410	0
	 ("00000000000000000000000000000000"),	 -- 1409	0
	 ("00000000000000000000000000000000"),	 -- 1408	0
	 ("00000000000000000000000000000000"),	 -- 1407	0
	 ("00000000000000000000000000000000"),	 -- 1406	0
	 ("00000000000000000000000000000000"),	 -- 1405	0
	 ("00000000000000000000000000000000"),	 -- 1404	0
	 ("00000000000000000000000000000000"),	 -- 1403	0
	 ("00000000000000000000000000000000"),	 -- 1402	0
	 ("00000000000000000000000000000000"),	 -- 1401	0
	 ("00000000000000000000000000000000"),	 -- 1400	0
	 ("00000000000000000000000000000000"),	 -- 1399	0
	 ("00000000000000000000000000000000"),	 -- 1398	0
	 ("00000000000000000000000000000000"),	 -- 1397	0
	 ("00000000000000000000000000000000"),	 -- 1396	0
	 ("00000000000000000000000000000000"),	 -- 1395	0
	 ("00000000000000000000000000000000"),	 -- 1394	0
	 ("00000000000000000000000000000000"),	 -- 1393	0
	 ("00000000000000000000000000000000"),	 -- 1392	0
	 ("00000000000000000000000000000000"),	 -- 1391	0
	 ("00000000000000000000000000000000"),	 -- 1390	0
	 ("00000000000000000000000000000000"),	 -- 1389	0
	 ("00000000000000000000000000000000"),	 -- 1388	0
	 ("00000000000000000000000000000000"),	 -- 1387	0
	 ("00000000000000000000000000000000"),	 -- 1386	0
	 ("00000000000000000000000000000000"),	 -- 1385	0
	 ("00000000000000000000000000000000"),	 -- 1384	0
	 ("00000000000000000000000000000000"),	 -- 1383	0
	 ("00000000000000000000000000000000"),	 -- 1382	0
	 ("00000000000000000000000000000000"),	 -- 1381	0
	 ("00000000000000000000000000000000"),	 -- 1380	0
	 ("00000000000000000000000000000000"),	 -- 1379	0
	 ("00000000000000000000000000000000"),	 -- 1378	0
	 ("00000000000000000000000000000000"),	 -- 1377	0
	 ("00000000000000000000000000000000"),	 -- 1376	0
	 ("00000000000000000000000000000000"),	 -- 1375	0
	 ("00000000000000000000000000000000"),	 -- 1374	0
	 ("00000000000000000000000000000000"),	 -- 1373	0
	 ("00000000000000000000000000000000"),	 -- 1372	0
	 ("00000000000000000000000000000000"),	 -- 1371	0
	 ("00000000000000000000000000000000"),	 -- 1370	0
	 ("00000000000000000000000000000000"),	 -- 1369	0
	 ("00000000000000000000000000000000"),	 -- 1368	0
	 ("00000000000000000000000000000000"),	 -- 1367	0
	 ("00000000000000000000000000000000"),	 -- 1366	0
	 ("00000000000000000000000000000000"),	 -- 1365	0
	 ("00000000000000000000000000000000"),	 -- 1364	0
	 ("00000000000000000000000000000000"),	 -- 1363	0
	 ("00000000000000000000000000000000"),	 -- 1362	0
	 ("00000000000000000000000000000000"),	 -- 1361	0
	 ("00000000000000000000000000000000"),	 -- 1360	0
	 ("00000000000000000000000000000000"),	 -- 1359	0
	 ("00000000000000000000000000000000"),	 -- 1358	0
	 ("00000000000000000000000000000000"),	 -- 1357	0
	 ("00000000000000000000000000000000"),	 -- 1356	0
	 ("00000000000000000000000000000000"),	 -- 1355	0
	 ("00000000000000000000000000000000"),	 -- 1354	0
	 ("00000000000000000000000000000000"),	 -- 1353	0
	 ("00000000000000000000000000000000"),	 -- 1352	0
	 ("00000000000000000000000000000000"),	 -- 1351	0
	 ("00000000000000000000000000000000"),	 -- 1350	0
	 ("00000000000000000000000000000000"),	 -- 1349	0
	 ("00000000000000000000000000000000"),	 -- 1348	0
	 ("00000000000000000000000000000000"),	 -- 1347	0
	 ("00000000000000000000000000000000"),	 -- 1346	0
	 ("00000000000000000000000000000000"),	 -- 1345	0
	 ("00000000000000000000000000000000"),	 -- 1344	0
	 ("00000000000000000000000000000000"),	 -- 1343	0
	 ("00000000000000000000000000000000"),	 -- 1342	0
	 ("00000000000000000000000000000000"),	 -- 1341	0
	 ("00000000000000000000000000000000"),	 -- 1340	0
	 ("00000000000000000000000000000000"),	 -- 1339	0
	 ("00000000000000000000000000000000"),	 -- 1338	0
	 ("00000000000000000000000000000000"),	 -- 1337	0
	 ("00000000000000000000000000000000"),	 -- 1336	0
	 ("00000000000000000000000000000000"),	 -- 1335	0
	 ("00000000000000000000000000000000"),	 -- 1334	0
	 ("00000000000000000000000000000000"),	 -- 1333	0
	 ("00000000000000000000000000000000"),	 -- 1332	0
	 ("00000000000000000000000000000000"),	 -- 1331	0
	 ("00000000000000000000000000000000"),	 -- 1330	0
	 ("00000000000000000000000000000000"),	 -- 1329	0
	 ("00000000000000000000000000000000"),	 -- 1328	0
	 ("00000000000000000000000000000000"),	 -- 1327	0
	 ("00000000000000000000000000000000"),	 -- 1326	0
	 ("00000000000000000000000000000000"),	 -- 1325	0
	 ("00000000000000000000000000000000"),	 -- 1324	0
	 ("00000000000000000000000000000000"),	 -- 1323	0
	 ("00000000000000000000000000000000"),	 -- 1322	0
	 ("00000000000000000000000000000000"),	 -- 1321	0
	 ("00000000000000000000000000000000"),	 -- 1320	0
	 ("00000000000000000000000000000000"),	 -- 1319	0
	 ("00000000000000000000000000000000"),	 -- 1318	0
	 ("00000000000000000000000000000000"),	 -- 1317	0
	 ("00000000000000000000000000000000"),	 -- 1316	0
	 ("00000000000000000000000000000000"),	 -- 1315	0
	 ("00000000000000000000000000000000"),	 -- 1314	0
	 ("00000000000000000000000000000000"),	 -- 1313	0
	 ("00000000000000000000000000000000"),	 -- 1312	0
	 ("00000000000000000000000000000000"),	 -- 1311	0
	 ("00000000000000000000000000000000"),	 -- 1310	0
	 ("00000000000000000000000000000000"),	 -- 1309	0
	 ("00000000000000000000000000000000"),	 -- 1308	0
	 ("00000000000000000000000000000000"),	 -- 1307	0
	 ("00000000000000000000000000000000"),	 -- 1306	0
	 ("00000000000000000000000000000000"),	 -- 1305	0
	 ("00000000000000000000000000000000"),	 -- 1304	0
	 ("00000000000000000000000000000000"),	 -- 1303	0
	 ("00000000000000000000000000000000"),	 -- 1302	0
	 ("00000000000000000000000000000000"),	 -- 1301	0
	 ("00000000000000000000000000000000"),	 -- 1300	0
	 ("00000000000000000000000000000000"),	 -- 1299	0
	 ("00000000000000000000000000000000"),	 -- 1298	0
	 ("00000000000000000000000000000000"),	 -- 1297	0
	 ("00000000000000000000000000000000"),	 -- 1296	0
	 ("00000000000000000000000000000000"),	 -- 1295	0
	 ("00000000000000000000000000000000"),	 -- 1294	0
	 ("00000000000000000000000000000000"),	 -- 1293	0
	 ("00000000000000000000000000000000"),	 -- 1292	0
	 ("00000000000000000000000000000000"),	 -- 1291	0
	 ("00000000000000000000000000000000"),	 -- 1290	0
	 ("00000000000000000000000000000000"),	 -- 1289	0
	 ("00000000000000000000000000000000"),	 -- 1288	0
	 ("00000000000000000000000000000000"),	 -- 1287	0
	 ("00000000000000000000000000000000"),	 -- 1286	0
	 ("00000000000000000000000000000000"),	 -- 1285	0
	 ("00000000000000000000000000000000"),	 -- 1284	0
	 ("00000000000000000000000000000000"),	 -- 1283	0
	 ("00000000000000000000000000000000"),	 -- 1282	0
	 ("00000000000000000000000000000000"),	 -- 1281	0
	 ("00000000000000000000000000000000"),	 -- 1280	0
	 ("00000000000000000000000000000000"),	 -- 1279	0
	 ("00000000000000000000000000000000"),	 -- 1278	0
	 ("00000000000000000000000000000000"),	 -- 1277	0
	 ("00000000000000000000000000000000"),	 -- 1276	0
	 ("00000000000000000000000000000000"),	 -- 1275	0
	 ("00000000000000000000000000000000"),	 -- 1274	0
	 ("00000000000000000000000000000000"),	 -- 1273	0
	 ("00000000000000000000000000000000"),	 -- 1272	0
	 ("00000000000000000000000000000000"),	 -- 1271	0
	 ("00000000000000000000000000000000"),	 -- 1270	0
	 ("00000000000000000000000000000000"),	 -- 1269	0
	 ("00000000000000000000000000000000"),	 -- 1268	0
	 ("00000000000000000000000000000000"),	 -- 1267	0
	 ("00000000000000000000000000000000"),	 -- 1266	0
	 ("00000000000000000000000000000000"),	 -- 1265	0
	 ("00000000000000000000000000000000"),	 -- 1264	0
	 ("00000000000000000000000000000000"),	 -- 1263	0
	 ("00000000000000000000000000000000"),	 -- 1262	0
	 ("00000000000000000000000000000000"),	 -- 1261	0
	 ("00000000000000000000000000000000"),	 -- 1260	0
	 ("00000000000000000000000000000000"),	 -- 1259	0
	 ("00000000000000000000000000000000"),	 -- 1258	0
	 ("00000000000000000000000000000000"),	 -- 1257	0
	 ("00000000000000000000000000000000"),	 -- 1256	0
	 ("00000000000000000000000000000000"),	 -- 1255	0
	 ("00000000000000000000000000000000"),	 -- 1254	0
	 ("00000000000000000000000000000000"),	 -- 1253	0
	 ("00000000000000000000000000000000"),	 -- 1252	0
	 ("00000000000000000000000000000000"),	 -- 1251	0
	 ("00000000000000000000000000000000"),	 -- 1250	0
	 ("00000000000000000000000000000000"),	 -- 1249	0
	 ("00000000000000000000000000000000"),	 -- 1248	0
	 ("00000000000000000000000000000000"),	 -- 1247	0
	 ("00000000000000000000000000000000"),	 -- 1246	0
	 ("00000000000000000000000000000000"),	 -- 1245	0
	 ("00000000000000000000000000000000"),	 -- 1244	0
	 ("00000000000000000000000000000000"),	 -- 1243	0
	 ("00000000000000000000000000000000"),	 -- 1242	0
	 ("00000000000000000000000000000000"),	 -- 1241	0
	 ("00000000000000000000000000000000"),	 -- 1240	0
	 ("00000000000000000000000000000000"),	 -- 1239	0
	 ("00000000000000000000000000000000"),	 -- 1238	0
	 ("00000000000000000000000000000000"),	 -- 1237	0
	 ("00000000000000000000000000000000"),	 -- 1236	0
	 ("00000000000000000000000000000000"),	 -- 1235	0
	 ("00000000000000000000000000000000"),	 -- 1234	0
	 ("00000000000000000000000000000000"),	 -- 1233	0
	 ("00000000000000000000000000000000"),	 -- 1232	0
	 ("00000000000000000000000000000000"),	 -- 1231	0
	 ("00000000000000000000000000000000"),	 -- 1230	0
	 ("00000000000000000000000000000000"),	 -- 1229	0
	 ("00000000000000000000000000000000"),	 -- 1228	0
	 ("00000000000000000000000000000000"),	 -- 1227	0
	 ("00000000000000000000000000000000"),	 -- 1226	0
	 ("00000000000000000000000000000000"),	 -- 1225	0
	 ("00000000000000000000000000000000"),	 -- 1224	0
	 ("00000000000000000000000000000000"),	 -- 1223	0
	 ("00000000000000000000000000000000"),	 -- 1222	0
	 ("00000000000000000000000000000000"),	 -- 1221	0
	 ("00000000000000000000000000000000"),	 -- 1220	0
	 ("00000000000000000000000000000000"),	 -- 1219	0
	 ("00000000000000000000000000000000"),	 -- 1218	0
	 ("00000000000000000000000000000000"),	 -- 1217	0
	 ("00000000000000000000000000000000"),	 -- 1216	0
	 ("00000000000000000000000000000000"),	 -- 1215	0
	 ("00000000000000000000000000000000"),	 -- 1214	0
	 ("00000000000000000000000000000000"),	 -- 1213	0
	 ("00000000000000000000000000000000"),	 -- 1212	0
	 ("00000000000000000000000000000000"),	 -- 1211	0
	 ("00000000000000000000000000000000"),	 -- 1210	0
	 ("00000000000000000000000000000000"),	 -- 1209	0
	 ("00000000000000000000000000000000"),	 -- 1208	0
	 ("00000000000000000000000000000000"),	 -- 1207	0
	 ("00000000000000000000000000000000"),	 -- 1206	0
	 ("00000000000000000000000000000000"),	 -- 1205	0
	 ("00000000000000000000000000000000"),	 -- 1204	0
	 ("00000000000000000000000000000000"),	 -- 1203	0
	 ("00000000000000000000000000000000"),	 -- 1202	0
	 ("00000000000000000000000000000000"),	 -- 1201	0
	 ("00000000000000000000000000000000"),	 -- 1200	0
	 ("00000000000000000000000000000000"),	 -- 1199	0
	 ("00000000000000000000000000000000"),	 -- 1198	0
	 ("00000000000000000000000000000000"),	 -- 1197	0
	 ("00000000000000000000000000000000"),	 -- 1196	0
	 ("00000000000000000000000000000000"),	 -- 1195	0
	 ("00000000000000000000000000000000"),	 -- 1194	0
	 ("00000000000000000000000000000000"),	 -- 1193	0
	 ("00000000000000000000000000000000"),	 -- 1192	0
	 ("00000000000000000000000000000000"),	 -- 1191	0
	 ("00000000000000000000000000000000"),	 -- 1190	0
	 ("00000000000000000000000000000000"),	 -- 1189	0
	 ("00000000000000000000000000000000"),	 -- 1188	0
	 ("00000000000000000000000000000000"),	 -- 1187	0
	 ("00000000000000000000000000000000"),	 -- 1186	0
	 ("00000000000000000000000000000000"),	 -- 1185	0
	 ("00000000000000000000000000000000"),	 -- 1184	0
	 ("00000000000000000000000000000000"),	 -- 1183	0
	 ("00000000000000000000000000000000"),	 -- 1182	0
	 ("00000000000000000000000000000000"),	 -- 1181	0
	 ("00000000000000000000000000000000"),	 -- 1180	0
	 ("00000000000000000000000000000000"),	 -- 1179	0
	 ("00000000000000000000000000000000"),	 -- 1178	0
	 ("00000000000000000000000000000000"),	 -- 1177	0
	 ("00000000000000000000000000000000"),	 -- 1176	0
	 ("00000000000000000000000000000000"),	 -- 1175	0
	 ("00000000000000000000000000000000"),	 -- 1174	0
	 ("00000000000000000000000000000000"),	 -- 1173	0
	 ("00000000000000000000000000000000"),	 -- 1172	0
	 ("00000000000000000000000000000000"),	 -- 1171	0
	 ("00000000000000000000000000000000"),	 -- 1170	0
	 ("00000000000000000000000000000000"),	 -- 1169	0
	 ("00000000000000000000000000000000"),	 -- 1168	0
	 ("00000000000000000000000000000000"),	 -- 1167	0
	 ("00000000000000000000000000000000"),	 -- 1166	0
	 ("00000000000000000000000000000000"),	 -- 1165	0
	 ("00000000000000000000000000000000"),	 -- 1164	0
	 ("00000000000000000000000000000000"),	 -- 1163	0
	 ("00000000000000000000000000000000"),	 -- 1162	0
	 ("00000000000000000000000000000000"),	 -- 1161	0
	 ("00000000000000000000000000000000"),	 -- 1160	0
	 ("00000000000000000000000000000000"),	 -- 1159	0
	 ("00000000000000000000000000000000"),	 -- 1158	0
	 ("00000000000000000000000000000000"),	 -- 1157	0
	 ("00000000000000000000000000000000"),	 -- 1156	0
	 ("00000000000000000000000000000000"),	 -- 1155	0
	 ("00000000000000000000000000000000"),	 -- 1154	0
	 ("00000000000000000000000000000000"),	 -- 1153	0
	 ("00000000000000000000000000000000"),	 -- 1152	0
	 ("00000000000000000000000000000000"),	 -- 1151	0
	 ("00000000000000000000000000000000"),	 -- 1150	0
	 ("00000000000000000000000000000000"),	 -- 1149	0
	 ("00000000000000000000000000000000"),	 -- 1148	0
	 ("00000000000000000000000000000000"),	 -- 1147	0
	 ("00000000000000000000000000000000"),	 -- 1146	0
	 ("00000000000000000000000000000000"),	 -- 1145	0
	 ("00000000000000000000000000000000"),	 -- 1144	0
	 ("00000000000000000000000000000000"),	 -- 1143	0
	 ("00000000000000000000000000000000"),	 -- 1142	0
	 ("00000000000000000000000000000000"),	 -- 1141	0
	 ("00000000000000000000000000000000"),	 -- 1140	0
	 ("00000000000000000000000000000000"),	 -- 1139	0
	 ("00000000000000000000000000000000"),	 -- 1138	0
	 ("00000000000000000000000000000000"),	 -- 1137	0
	 ("00000000000000000000000000000000"),	 -- 1136	0
	 ("00000000000000000000000000000000"),	 -- 1135	0
	 ("00000000000000000000000000000000"),	 -- 1134	0
	 ("00000000000000000000000000000000"),	 -- 1133	0
	 ("00000000000000000000000000000000"),	 -- 1132	0
	 ("00000000000000000000000000000000"),	 -- 1131	0
	 ("00000000000000000000000000000000"),	 -- 1130	0
	 ("00000000000000000000000000000000"),	 -- 1129	0
	 ("00000000000000000000000000000000"),	 -- 1128	0
	 ("00000000000000000000000000000000"),	 -- 1127	0
	 ("00000000000000000000000000000000"),	 -- 1126	0
	 ("00000000000000000000000000000000"),	 -- 1125	0
	 ("00000000000000000000000000000000"),	 -- 1124	0
	 ("00000000000000000000000000000000"),	 -- 1123	0
	 ("00000000000000000000000000000000"),	 -- 1122	0
	 ("00000000000000000000000000000000"),	 -- 1121	0
	 ("00000000000000000000000000000000"),	 -- 1120	0
	 ("00000000000000000000000000000000"),	 -- 1119	0
	 ("00000000000000000000000000000000"),	 -- 1118	0
	 ("00000000000000000000000000000000"),	 -- 1117	0
	 ("00000000000000000000000000000000"),	 -- 1116	0
	 ("00000000000000000000000000000000"),	 -- 1115	0
	 ("00000000000000000000000000000000"),	 -- 1114	0
	 ("00000000000000000000000000000000"),	 -- 1113	0
	 ("00000000000000000000000000000000"),	 -- 1112	0
	 ("00000000000000000000000000000000"),	 -- 1111	0
	 ("00000000000000000000000000000000"),	 -- 1110	0
	 ("00000000000000000000000000000000"),	 -- 1109	0
	 ("00000000000000000000000000000000"),	 -- 1108	0
	 ("00000000000000000000000000000000"),	 -- 1107	0
	 ("00000000000000000000000000000000"),	 -- 1106	0
	 ("00000000000000000000000000000000"),	 -- 1105	0
	 ("00000000000000000000000000000000"),	 -- 1104	0
	 ("00000000000000000000000000000000"),	 -- 1103	0
	 ("00000000000000000000000000000000"),	 -- 1102	0
	 ("00000000000000000000000000000000"),	 -- 1101	0
	 ("00000000000000000000000000000000"),	 -- 1100	0
	 ("00000000000000000000000000000000"),	 -- 1099	0
	 ("00000000000000000000000000000000"),	 -- 1098	0
	 ("00000000000000000000000000000000"),	 -- 1097	0
	 ("00000000000000000000000000000000"),	 -- 1096	0
	 ("00000000000000000000000000000000"),	 -- 1095	0
	 ("00000000000000000000000000000000"),	 -- 1094	0
	 ("00000000000000000000000000000000"),	 -- 1093	0
	 ("00000000000000000000000000000000"),	 -- 1092	0
	 ("00000000000000000000000000000000"),	 -- 1091	0
	 ("00000000000000000000000000000000"),	 -- 1090	0
	 ("00000000000000000000000000000000"),	 -- 1089	0
	 ("00000000000000000000000000000000"),	 -- 1088	0
	 ("00000000000000000000000000000000"),	 -- 1087	0
	 ("00000000000000000000000000000000"),	 -- 1086	0
	 ("00000000000000000000000000000000"),	 -- 1085	0
	 ("00000000000000000000000000000000"),	 -- 1084	0
	 ("00000000000000000000000000000000"),	 -- 1083	0
	 ("00000000000000000000000000000000"),	 -- 1082	0
	 ("00000000000000000000000000000000"),	 -- 1081	0
	 ("00000000000000000000000000000000"),	 -- 1080	0
	 ("00000000000000000000000000000000"),	 -- 1079	0
	 ("00000000000000000000000000000000"),	 -- 1078	0
	 ("00000000000000000000000000000000"),	 -- 1077	0
	 ("00000000000000000000000000000000"),	 -- 1076	0
	 ("00000000000000000000000000000000"),	 -- 1075	0
	 ("00000000000000000000000000000000"),	 -- 1074	0
	 ("00000000000000000000000000000000"),	 -- 1073	0
	 ("00000000000000000000000000000000"),	 -- 1072	0
	 ("00000000000000000000000000000000"),	 -- 1071	0
	 ("00000000000000000000000000000000"),	 -- 1070	0
	 ("00000000000000000000000000000000"),	 -- 1069	0
	 ("00000000000000000000000000000000"),	 -- 1068	0
	 ("00000000000000000000000000000000"),	 -- 1067	0
	 ("00000000000000000000000000000000"),	 -- 1066	0
	 ("00000000000000000000000000000000"),	 -- 1065	0
	 ("00000000000000000000000000000000"),	 -- 1064	0
	 ("00000000000000000000000000000000"),	 -- 1063	0
	 ("00000000000000000000000000000000"),	 -- 1062	0
	 ("00000000000000000000000000000000"),	 -- 1061	0
	 ("00000000000000000000000000000000"),	 -- 1060	0
	 ("00000000000000000000000000000000"),	 -- 1059	0
	 ("00000000000000000000000000000000"),	 -- 1058	0
	 ("00000000000000000000000000000000"),	 -- 1057	0
	 ("00000000000000000000000000000000"),	 -- 1056	0
	 ("00000000000000000000000000000000"),	 -- 1055	0
	 ("00000000000000000000000000000000"),	 -- 1054	0
	 ("00000000000000000000000000000000"),	 -- 1053	0
	 ("00000000000000000000000000000000"),	 -- 1052	0
	 ("00000000000000000000000000000000"),	 -- 1051	0
	 ("00000000000000000000000000000000"),	 -- 1050	0
	 ("00000000000000000000000000000000"),	 -- 1049	0
	 ("00000000000000000000000000000000"),	 -- 1048	0
	 ("00000000000000000000000000000000"),	 -- 1047	0
	 ("00000000000000000000000000000000"),	 -- 1046	0
	 ("00000000000000000000000000000000"),	 -- 1045	0
	 ("00000000000000000000000000000000"),	 -- 1044	0
	 ("00000000000000000000000000000000"),	 -- 1043	0
	 ("00000000000000000000000000000000"),	 -- 1042	0
	 ("00000000000000000000000000000000"),	 -- 1041	0
	 ("00000000000000000000000000000000"),	 -- 1040	0
	 ("00000000000000000000000000000000"),	 -- 1039	0
	 ("00000000000000000000000000000000"),	 -- 1038	0
	 ("00000000000000000000000000000000"),	 -- 1037	0
	 ("00000000000000000000000000000000"),	 -- 1036	0
	 ("00000000000000000000000000000000"),	 -- 1035	0
	 ("00000000000000000000000000000000"),	 -- 1034	0
	 ("00000000000000000000000000000000"),	 -- 1033	0
	 ("00000000000000000000000000000000"),	 -- 1032	0
	 ("00000000000000000000000000000000"),	 -- 1031	0
	 ("00000000000000000000000000000000"),	 -- 1030	0
	 ("00000000000000000000000000000000"),	 -- 1029	0
	 ("00000000000000000000000000000000"),	 -- 1028	0
	 ("00000000000000000000000000000000"),	 -- 1027	0
	 ("00000000000000000000000000000000"),	 -- 1026	0
	 ("00000000000000000000000000000000"),	 -- 1025	0
	 ("00000000000000000000000000000000"),	 -- 1024	0
	 ("00000000000000000000000000000000"),	 -- 1023	0
	 ("00000000000000000000000000000000"),	 -- 1022	0
	 ("00000000000000000000000000000000"),	 -- 1021	0
	 ("00000000000000000000000000000000"),	 -- 1020	0
	 ("00000000000000000000000000000000"),	 -- 1019	0
	 ("00000000000000000000000000000000"),	 -- 1018	0
	 ("00000000000000000000000000000000"),	 -- 1017	0
	 ("00000000000000000000000000000000"),	 -- 1016	0
	 ("00000000000000000000000000000000"),	 -- 1015	0
	 ("00000000000000000000000000000000"),	 -- 1014	0
	 ("00000000000000000000000000000000"),	 -- 1013	0
	 ("00000000000000000000000000000000"),	 -- 1012	0
	 ("00000000000000000000000000000000"),	 -- 1011	0
	 ("00000000000000000000000000000000"),	 -- 1010	0
	 ("00000000000000000000000000000000"),	 -- 1009	0
	 ("00000000000000000000000000000000"),	 -- 1008	0
	 ("00000000000000000000000000000000"),	 -- 1007	0
	 ("00000000000000000000000000000000"),	 -- 1006	0
	 ("00000000000000000000000000000000"),	 -- 1005	0
	 ("00000000000000000000000000000000"),	 -- 1004	0
	 ("00000000000000000000000000000000"),	 -- 1003	0
	 ("00000000000000000000000000000000"),	 -- 1002	0
	 ("00000000000000000000000000000000"),	 -- 1001	0
	 ("00000000000000000000000000000000"),	 -- 1000	0
	 ("00000000000000000000000000000000"),	 -- 999	0
	 ("00000000000000000000000000000000"),	 -- 998	0
	 ("00000000000000000000000000000000"),	 -- 997	0
	 ("00000000000000000000000000000000"),	 -- 996	0
	 ("00000000000000000000000000000000"),	 -- 995	0
	 ("00000000000000000000000000000000"),	 -- 994	0
	 ("00000000000000000000000000000000"),	 -- 993	0
	 ("00000000000000000000000000000000"),	 -- 992	0
	 ("00000000000000000000000000000000"),	 -- 991	0
	 ("00000000000000000000000000000000"),	 -- 990	0
	 ("00000000000000000000000000000000"),	 -- 989	0
	 ("00000000000000000000000000000000"),	 -- 988	0
	 ("00000000000000000000000000000000"),	 -- 987	0
	 ("00000000000000000000000000000000"),	 -- 986	0
	 ("00000000000000000000000000000000"),	 -- 985	0
	 ("00000000000000000000000000000000"),	 -- 984	0
	 ("00000000000000000000000000000000"),	 -- 983	0
	 ("00000000000000000000000000000000"),	 -- 982	0
	 ("00000000000000000000000000000000"),	 -- 981	0
	 ("00000000000000000000000000000000"),	 -- 980	0
	 ("00000000000000000000000000000000"),	 -- 979	0
	 ("00000000000000000000000000000000"),	 -- 978	0
	 ("00000000000000000000000000000000"),	 -- 977	0
	 ("00000000000000000000000000000000"),	 -- 976	0
	 ("00000000000000000000000000000000"),	 -- 975	0
	 ("00000000000000000000000000000000"),	 -- 974	0
	 ("00000000000000000000000000000000"),	 -- 973	0
	 ("00000000000000000000000000000000"),	 -- 972	0
	 ("00000000000000000000000000000000"),	 -- 971	0
	 ("00000000000000000000000000000000"),	 -- 970	0
	 ("00000000000000000000000000000000"),	 -- 969	0
	 ("00000000000000000000000000000000"),	 -- 968	0
	 ("00000000000000000000000000000000"),	 -- 967	0
	 ("00000000000000000000000000000000"),	 -- 966	0
	 ("00000000000000000000000000000000"),	 -- 965	0
	 ("00000000000000000000000000000000"),	 -- 964	0
	 ("00000000000000000000000000000000"),	 -- 963	0
	 ("00000000000000000000000000000000"),	 -- 962	0
	 ("00000000000000000000000000000000"),	 -- 961	0
	 ("00000000000000000000000000000000"),	 -- 960	0
	 ("00000000000000000000000000000000"),	 -- 959	0
	 ("00000000000000000000000000000000"),	 -- 958	0
	 ("00000000000000000000000000000000"),	 -- 957	0
	 ("00000000000000000000000000000000"),	 -- 956	0
	 ("00000000000000000000000000000000"),	 -- 955	0
	 ("00000000000000000000000000000000"),	 -- 954	0
	 ("00000000000000000000000000000000"),	 -- 953	0
	 ("00000000000000000000000000000000"),	 -- 952	0
	 ("00000000000000000000000000000000"),	 -- 951	0
	 ("00000000000000000000000000000000"),	 -- 950	0
	 ("00000000000000000000000000000000"),	 -- 949	0
	 ("00000000000000000000000000000000"),	 -- 948	0
	 ("00000000000000000000000000000000"),	 -- 947	0
	 ("00000000000000000000000000000000"),	 -- 946	0
	 ("00000000000000000000000000000000"),	 -- 945	0
	 ("00000000000000000000000000000000"),	 -- 944	0
	 ("00000000000000000000000000000000"),	 -- 943	0
	 ("00000000000000000000000000000000"),	 -- 942	0
	 ("00000000000000000000000000000000"),	 -- 941	0
	 ("00000000000000000000000000000000"),	 -- 940	0
	 ("00000000000000000000000000000000"),	 -- 939	0
	 ("00000000000000000000000000000000"),	 -- 938	0
	 ("00000000000000000000000000000000"),	 -- 937	0
	 ("00000000000000000000000000000000"),	 -- 936	0
	 ("00000000000000000000000000000000"),	 -- 935	0
	 ("00000000000000000000000000000000"),	 -- 934	0
	 ("00000000000000000000000000000000"),	 -- 933	0
	 ("00000000000000000000000000000000"),	 -- 932	0
	 ("00000000000000000000000000000000"),	 -- 931	0
	 ("00000000000000000000000000000000"),	 -- 930	0
	 ("00000000000000000000000000000000"),	 -- 929	0
	 ("00000000000000000000000000000000"),	 -- 928	0
	 ("00000000000000000000000000000000"),	 -- 927	0
	 ("00000000000000000000000000000000"),	 -- 926	0
	 ("00000000000000000000000000000000"),	 -- 925	0
	 ("00000000000000000000000000000000"),	 -- 924	0
	 ("00000000000000000000000000000000"),	 -- 923	0
	 ("00000000000000000000000000000000"),	 -- 922	0
	 ("00000000000000000000000000000000"),	 -- 921	0
	 ("00000000000000000000000000000000"),	 -- 920	0
	 ("00000000000000000000000000000000"),	 -- 919	0
	 ("00000000000000000000000000000000"),	 -- 918	0
	 ("00000000000000000000000000000000"),	 -- 917	0
	 ("00000000000000000000000000000000"),	 -- 916	0
	 ("00000000000000000000000000000000"),	 -- 915	0
	 ("00000000000000000000000000000000"),	 -- 914	0
	 ("00000000000000000000000000000000"),	 -- 913	0
	 ("00000000000000000000000000000000"),	 -- 912	0
	 ("00000000000000000000000000000000"),	 -- 911	0
	 ("00000000000000000000000000000000"),	 -- 910	0
	 ("00000000000000000000000000000000"),	 -- 909	0
	 ("00000000000000000000000000000000"),	 -- 908	0
	 ("00000000000000000000000000000000"),	 -- 907	0
	 ("00000000000000000000000000000000"),	 -- 906	0
	 ("00000000000000000000000000000000"),	 -- 905	0
	 ("00000000000000000000000000000000"),	 -- 904	0
	 ("00000000000000000000000000000000"),	 -- 903	0
	 ("00000000000000000000000000000000"),	 -- 902	0
	 ("00000000000000000000000000000000"),	 -- 901	0
	 ("00000000000000000000000000000000"),	 -- 900	0
	 ("00000000000000000000000000000000"),	 -- 899	0
	 ("00000000000000000000000000000000"),	 -- 898	0
	 ("00000000000000000000000000000000"),	 -- 897	0
	 ("00000000000000000000000000000000"),	 -- 896	0
	 ("00000000000000000000000000000000"),	 -- 895	0
	 ("00000000000000000000000000000000"),	 -- 894	0
	 ("00000000000000000000000000000000"),	 -- 893	0
	 ("00000000000000000000000000000000"),	 -- 892	0
	 ("00000000000000000000000000000000"),	 -- 891	0
	 ("00000000000000000000000000000000"),	 -- 890	0
	 ("00000000000000000000000000000000"),	 -- 889	0
	 ("00000000000000000000000000000000"),	 -- 888	0
	 ("00000000000000000000000000000000"),	 -- 887	0
	 ("00000000000000000000000000000000"),	 -- 886	0
	 ("00000000000000000000000000000000"),	 -- 885	0
	 ("00000000000000000000000000000000"),	 -- 884	0
	 ("00000000000000000000000000000000"),	 -- 883	0
	 ("00000000000000000000000000000000"),	 -- 882	0
	 ("00000000000000000000000000000000"),	 -- 881	0
	 ("00000000000000000000000000000000"),	 -- 880	0
	 ("00000000000000000000000000000000"),	 -- 879	0
	 ("00000000000000000000000000000000"),	 -- 878	0
	 ("00000000000000000000000000000000"),	 -- 877	0
	 ("00000000000000000000000000000000"),	 -- 876	0
	 ("00000000000000000000000000000000"),	 -- 875	0
	 ("00000000000000000000000000000000"),	 -- 874	0
	 ("00000000000000000000000000000000"),	 -- 873	0
	 ("00000000000000000000000000000000"),	 -- 872	0
	 ("00000000000000000000000000000000"),	 -- 871	0
	 ("00000000000000000000000000000000"),	 -- 870	0
	 ("00000000000000000000000000000000"),	 -- 869	0
	 ("00000000000000000000000000000000"),	 -- 868	0
	 ("00000000000000000000000000000000"),	 -- 867	0
	 ("00000000000000000000000000000000"),	 -- 866	0
	 ("00000000000000000000000000000000"),	 -- 865	0
	 ("00000000000000000000000000000000"),	 -- 864	0
	 ("00000000000000000000000000000000"),	 -- 863	0
	 ("00000000000000000000000000000000"),	 -- 862	0
	 ("00000000000000000000000000000000"),	 -- 861	0
	 ("00000000000000000000000000000000"),	 -- 860	0
	 ("00000000000000000000000000000000"),	 -- 859	0
	 ("00000000000000000000000000000000"),	 -- 858	0
	 ("00000000000000000000000000000000"),	 -- 857	0
	 ("00000000000000000000000000000000"),	 -- 856	0
	 ("00000000000000000000000000000000"),	 -- 855	0
	 ("00000000000000000000000000000000"),	 -- 854	0
	 ("00000000000000000000000000000000"),	 -- 853	0
	 ("00000000000000000000000000000000"),	 -- 852	0
	 ("00000000000000000000000000000000"),	 -- 851	0
	 ("00000000000000000000000000000000"),	 -- 850	0
	 ("00000000000000000000000000000000"),	 -- 849	0
	 ("00000000000000000000000000000000"),	 -- 848	0
	 ("00000000000000000000000000000000"),	 -- 847	0
	 ("00000000000000000000000000000000"),	 -- 846	0
	 ("00000000000000000000000000000000"),	 -- 845	0
	 ("00000000000000000000000000000000"),	 -- 844	0
	 ("00000000000000000000000000000000"),	 -- 843	0
	 ("00000000000000000000000000000000"),	 -- 842	0
	 ("00000000000000000000000000000000"),	 -- 841	0
	 ("00000000000000000000000000000000"),	 -- 840	0
	 ("00000000000000000000000000000000"),	 -- 839	0
	 ("00000000000000000000000000000000"),	 -- 838	0
	 ("00000000000000000000000000000000"),	 -- 837	0
	 ("00000000000000000000000000000000"),	 -- 836	0
	 ("00000000000000000000000000000000"),	 -- 835	0
	 ("00000000000000000000000000000000"),	 -- 834	0
	 ("00000000000000000000000000000000"),	 -- 833	0
	 ("00000000000000000000000000000000"),	 -- 832	0
	 ("00000000000000000000000000000000"),	 -- 831	0
	 ("00000000000000000000000000000000"),	 -- 830	0
	 ("00000000000000000000000000000000"),	 -- 829	0
	 ("00000000000000000000000000000000"),	 -- 828	0
	 ("00000000000000000000000000000000"),	 -- 827	0
	 ("00000000000000000000000000000000"),	 -- 826	0
	 ("00000000000000000000000000000000"),	 -- 825	0
	 ("00000000000000000000000000000000"),	 -- 824	0
	 ("00000000000000000000000000000000"),	 -- 823	0
	 ("00000000000000000000000000000000"),	 -- 822	0
	 ("00000000000000000000000000000000"),	 -- 821	0
	 ("00000000000000000000000000000000"),	 -- 820	0
	 ("00000000000000000000000000000000"),	 -- 819	0
	 ("00000000000000000000000000000000"),	 -- 818	0
	 ("00000000000000000000000000000000"),	 -- 817	0
	 ("00000000000000000000000000000000"),	 -- 816	0
	 ("00000000000000000000000000000000"),	 -- 815	0
	 ("00000000000000000000000000000000"),	 -- 814	0
	 ("00000000000000000000000000000000"),	 -- 813	0
	 ("00000000000000000000000000000000"),	 -- 812	0
	 ("00000000000000000000000000000000"),	 -- 811	0
	 ("00000000000000000000000000000000"),	 -- 810	0
	 ("00000000000000000000000000000000"),	 -- 809	0
	 ("00000000000000000000000000000000"),	 -- 808	0
	 ("00000000000000000000000000000000"),	 -- 807	0
	 ("00000000000000000000000000000000"),	 -- 806	0
	 ("00000000000000000000000000000000"),	 -- 805	0
	 ("00000000000000000000000000000000"),	 -- 804	0
	 ("00000000000000000000000000000000"),	 -- 803	0
	 ("00000000000000000000000000000000"),	 -- 802	0
	 ("00000000000000000000000000000000"),	 -- 801	0
	 ("00000000000000000000000000000000"),	 -- 800	0
	 ("00000000000000000000000000000000"),	 -- 799	0
	 ("00000000000000000000000000000000"),	 -- 798	0
	 ("00000000000000000000000000000000"),	 -- 797	0
	 ("00000000000000000000000000000000"),	 -- 796	0
	 ("00000000000000000000000000000000"),	 -- 795	0
	 ("00000000000000000000000000000000"),	 -- 794	0
	 ("00000000000000000000000000000000"),	 -- 793	0
	 ("00000000000000000000000000000000"),	 -- 792	0
	 ("00000000000000000000000000000000"),	 -- 791	0
	 ("00000000000000000000000000000000"),	 -- 790	0
	 ("00000000000000000000000000000000"),	 -- 789	0
	 ("00000000000000000000000000000000"),	 -- 788	0
	 ("00000000000000000000000000000000"),	 -- 787	0
	 ("00000000000000000000000000000000"),	 -- 786	0
	 ("00000000000000000000000000000000"),	 -- 785	0
	 ("00000000000000000000000000000000"),	 -- 784	0
	 ("00000000000000000000000000000000"),	 -- 783	0
	 ("00000000000000000000000000000000"),	 -- 782	0
	 ("00000000000000000000000000000000"),	 -- 781	0
	 ("00000000000000000000000000000000"),	 -- 780	0
	 ("00000000000000000000000000000000"),	 -- 779	0
	 ("00000000000000000000000000000000"),	 -- 778	0
	 ("00000000000000000000000000000000"),	 -- 777	0
	 ("00000000000000000000000000000000"),	 -- 776	0
	 ("00000000000000000000000000000000"),	 -- 775	0
	 ("00000000000000000000000000000000"),	 -- 774	0
	 ("00000000000000000000000000000000"),	 -- 773	0
	 ("00000000000000000000000000000000"),	 -- 772	0
	 ("00000000000000000000000000000000"),	 -- 771	0
	 ("00000000000000000000000000000000"),	 -- 770	0
	 ("00000000000000000000000000000000"),	 -- 769	0
	 ("00000000000000000000000000000000"),	 -- 768	0
	 ("00000000000000000000000000000000"),	 -- 767	0
	 ("00000000000000000000000000000000"),	 -- 766	0
	 ("00000000000000000000000000000000"),	 -- 765	0
	 ("00000000000000000000000000000000"),	 -- 764	0
	 ("00000000000000000000000000000000"),	 -- 763	0
	 ("00000000000000000000000000000000"),	 -- 762	0
	 ("00000000000000000000000000000000"),	 -- 761	0
	 ("00000000000000000000000000000000"),	 -- 760	0
	 ("00000000000000000000000000000000"),	 -- 759	0
	 ("00000000000000000000000000000000"),	 -- 758	0
	 ("00000000000000000000000000000000"),	 -- 757	0
	 ("00000000000000000000000000000000"),	 -- 756	0
	 ("00000000000000000000000000000000"),	 -- 755	0
	 ("00000000000000000000000000000000"),	 -- 754	0
	 ("00000000000000000000000000000000"),	 -- 753	0
	 ("00000000000000000000000000000000"),	 -- 752	0
	 ("00000000000000000000000000000000"),	 -- 751	0
	 ("00000000000000000000000000000000"),	 -- 750	0
	 ("00000000000000000000000000000000"),	 -- 749	0
	 ("00000000000000000000000000000000"),	 -- 748	0
	 ("00000000000000000000000000000000"),	 -- 747	0
	 ("00000000000000000000000000000000"),	 -- 746	0
	 ("00000000000000000000000000000000"),	 -- 745	0
	 ("00000000000000000000000000000000"),	 -- 744	0
	 ("00000000000000000000000000000000"),	 -- 743	0
	 ("00000000000000000000000000000000"),	 -- 742	0
	 ("00000000000000000000000000000000"),	 -- 741	0
	 ("00000000000000000000000000000000"),	 -- 740	0
	 ("00000000000000000000000000000000"),	 -- 739	0
	 ("00000000000000000000000000000000"),	 -- 738	0
	 ("00000000000000000000000000000000"),	 -- 737	0
	 ("00000000000000000000000000000000"),	 -- 736	0
	 ("00000000000000000000000000000000"),	 -- 735	0
	 ("00000000000000000000000000000000"),	 -- 734	0
	 ("00000000000000000000000000000000"),	 -- 733	0
	 ("00000000000000000000000000000000"),	 -- 732	0
	 ("00000000000000000000000000000000"),	 -- 731	0
	 ("00000000000000000000000000000000"),	 -- 730	0
	 ("00000000000000000000000000000000"),	 -- 729	0
	 ("00000000000000000000000000000000"),	 -- 728	0
	 ("00000000000000000000000000000000"),	 -- 727	0
	 ("00000000000000000000000000000000"),	 -- 726	0
	 ("00000000000000000000000000000000"),	 -- 725	0
	 ("00000000000000000000000000000000"),	 -- 724	0
	 ("00000000000000000000000000000000"),	 -- 723	0
	 ("00000000000000000000000000000000"),	 -- 722	0
	 ("00000000000000000000000000000000"),	 -- 721	0
	 ("00000000000000000000000000000000"),	 -- 720	0
	 ("00000000000000000000000000000000"),	 -- 719	0
	 ("00000000000000000000000000000000"),	 -- 718	0
	 ("00000000000000000000000000000000"),	 -- 717	0
	 ("00000000000000000000000000000000"),	 -- 716	0
	 ("00000000000000000000000000000000"),	 -- 715	0
	 ("00000000000000000000000000000000"),	 -- 714	0
	 ("00000000000000000000000000000000"),	 -- 713	0
	 ("00000000000000000000000000000000"),	 -- 712	0
	 ("00000000000000000000000000000000"),	 -- 711	0
	 ("00000000000000000000000000000000"),	 -- 710	0
	 ("00000000000000000000000000000000"),	 -- 709	0
	 ("00000000000000000000000000000000"),	 -- 708	0
	 ("00000000000000000000000000000000"),	 -- 707	0
	 ("00000000000000000000000000000000"),	 -- 706	0
	 ("00000000000000000000000000000000"),	 -- 705	0
	 ("00000000000000000000000000000000"),	 -- 704	0
	 ("00000000000000000000000000000000"),	 -- 703	0
	 ("00000000000000000000000000000000"),	 -- 702	0
	 ("00000000000000000000000000000000"),	 -- 701	0
	 ("00000000000000000000000000000000"),	 -- 700	0
	 ("00000000000000000000000000000000"),	 -- 699	0
	 ("00000000000000000000000000000000"),	 -- 698	0
	 ("00000000000000000000000000000000"),	 -- 697	0
	 ("00000000000000000000000000000000"),	 -- 696	0
	 ("00000000000000000000000000000000"),	 -- 695	0
	 ("00000000000000000000000000000000"),	 -- 694	0
	 ("00000000000000000000000000000000"),	 -- 693	0
	 ("00000000000000000000000000000000"),	 -- 692	0
	 ("00000000000000000000000000000000"),	 -- 691	0
	 ("00000000000000000000000000000000"),	 -- 690	0
	 ("00000000000000000000000000000000"),	 -- 689	0
	 ("00000000000000000000000000000000"),	 -- 688	0
	 ("00000000000000000000000000000000"),	 -- 687	0
	 ("00000000000000000000000000000000"),	 -- 686	0
	 ("00000000000000000000000000000000"),	 -- 685	0
	 ("00000000000000000000000000000000"),	 -- 684	0
	 ("00000000000000000000000000000000"),	 -- 683	0
	 ("00000000000000000000000000000000"),	 -- 682	0
	 ("00000000000000000000000000000000"),	 -- 681	0
	 ("00000000000000000000000000000000"),	 -- 680	0
	 ("00000000000000000000000000000000"),	 -- 679	0
	 ("00000000000000000000000000000000"),	 -- 678	0
	 ("00000000000000000000000000000000"),	 -- 677	0
	 ("00000000000000000000000000000000"),	 -- 676	0
	 ("00000000000000000000000000000000"),	 -- 675	0
	 ("00000000000000000000000000000000"),	 -- 674	0
	 ("00000000000000000000000000000000"),	 -- 673	0
	 ("00000000000000000000000000000000"),	 -- 672	0
	 ("00000000000000000000000000000000"),	 -- 671	0
	 ("00000000000000000000000000000000"),	 -- 670	0
	 ("00000000000000000000000000000000"),	 -- 669	0
	 ("00000000000000000000000000000000"),	 -- 668	0
	 ("00000000000000000000000000000000"),	 -- 667	0
	 ("00000000000000000000000000000000"),	 -- 666	0
	 ("00000000000000000000000000000000"),	 -- 665	0
	 ("00000000000000000000000000000000"),	 -- 664	0
	 ("00000000000000000000000000000000"),	 -- 663	0
	 ("00000000000000000000000000000000"),	 -- 662	0
	 ("00000000000000000000000000000000"),	 -- 661	0
	 ("00000000000000000000000000000000"),	 -- 660	0
	 ("00000000000000000000000000000000"),	 -- 659	0
	 ("00000000000000000000000000000000"),	 -- 658	0
	 ("00000000000000000000000000000000"),	 -- 657	0
	 ("00000000000000000000000000000000"),	 -- 656	0
	 ("00000000000000000000000000000000"),	 -- 655	0
	 ("00000000000000000000000000000000"),	 -- 654	0
	 ("00000000000000000000000000000000"),	 -- 653	0
	 ("00000000000000000000000000000000"),	 -- 652	0
	 ("00000000000000000000000000000000"),	 -- 651	0
	 ("00000000000000000000000000000000"),	 -- 650	0
	 ("00000000000000000000000000000000"),	 -- 649	0
	 ("00000000000000000000000000000000"),	 -- 648	0
	 ("00000000000000000000000000000000"),	 -- 647	0
	 ("00000000000000000000000000000000"),	 -- 646	0
	 ("00000000000000000000000000000000"),	 -- 645	0
	 ("00000000000000000000000000000000"),	 -- 644	0
	 ("00000000000000000000000000000000"),	 -- 643	0
	 ("00000000000000000000000000000000"),	 -- 642	0
	 ("00000000000000000000000000000000"),	 -- 641	0
	 ("00000000000000000000000000000000"),	 -- 640	0
	 ("00000000000000000000000000000000"),	 -- 639	0
	 ("00000000000000000000000000000000"),	 -- 638	0
	 ("00000000000000000000000000000000"),	 -- 637	0
	 ("00000000000000000000000000000000"),	 -- 636	0
	 ("00000000000000000000000000000000"),	 -- 635	0
	 ("00000000000000000000000000000000"),	 -- 634	0
	 ("00000000000000000000000000000000"),	 -- 633	0
	 ("00000000000000000000000000000000"),	 -- 632	0
	 ("00000000000000000000000000000000"),	 -- 631	0
	 ("00000000000000000000000000000000"),	 -- 630	0
	 ("00000000000000000000000000000000"),	 -- 629	0
	 ("00000000000000000000000000000000"),	 -- 628	0
	 ("00000000000000000000000000000000"),	 -- 627	0
	 ("00000000000000000000000000000000"),	 -- 626	0
	 ("00000000000000000000000000000000"),	 -- 625	0
	 ("00000000000000000000000000000000"),	 -- 624	0
	 ("00000000000000000000000000000000"),	 -- 623	0
	 ("00000000000000000000000000000000"),	 -- 622	0
	 ("00000000000000000000000000000000"),	 -- 621	0
	 ("00000000000000000000000000000000"),	 -- 620	0
	 ("00000000000000000000000000000000"),	 -- 619	0
	 ("00000000000000000000000000000000"),	 -- 618	0
	 ("00000000000000000000000000000000"),	 -- 617	0
	 ("00000000000000000000000000000000"),	 -- 616	0
	 ("00000000000000000000000000000000"),	 -- 615	0
	 ("00000000000000000000000000000000"),	 -- 614	0
	 ("00000000000000000000000000000000"),	 -- 613	0
	 ("00000000000000000000000000000000"),	 -- 612	0
	 ("00000000000000000000000000000000"),	 -- 611	0
	 ("00000000000000000000000000000000"),	 -- 610	0
	 ("00000000000000000000000000000000"),	 -- 609	0
	 ("00000000000000000000000000000000"),	 -- 608	0
	 ("00000000000000000000000000000000"),	 -- 607	0
	 ("00000000000000000000000000000000"),	 -- 606	0
	 ("00000000000000000000000000000000"),	 -- 605	0
	 ("00000000000000000000000000000000"),	 -- 604	0
	 ("00000000000000000000000000000000"),	 -- 603	0
	 ("00000000000000000000000000000000"),	 -- 602	0
	 ("00000000000000000000000000000000"),	 -- 601	0
	 ("00000000000000000000000000000000"),	 -- 600	0
	 ("00000000000000000000000000000000"),	 -- 599	0
	 ("00000000000000000000000000000000"),	 -- 598	0
	 ("00000000000000000000000000000000"),	 -- 597	0
	 ("00000000000000000000000000000000"),	 -- 596	0
	 ("00000000000000000000000000000000"),	 -- 595	0
	 ("00000000000000000000000000000000"),	 -- 594	0
	 ("00000000000000000000000000000000"),	 -- 593	0
	 ("00000000000000000000000000000000"),	 -- 592	0
	 ("00000000000000000000000000000000"),	 -- 591	0
	 ("00000000000000000000000000000000"),	 -- 590	0
	 ("00000000000000000000000000000000"),	 -- 589	0
	 ("00000000000000000000000000000000"),	 -- 588	0
	 ("00000000000000000000000000000000"),	 -- 587	0
	 ("00000000000000000000000000000000"),	 -- 586	0
	 ("00000000000000000000000000000000"),	 -- 585	0
	 ("00000000000000000000000000000000"),	 -- 584	0
	 ("00000000000000000000000000000000"),	 -- 583	0
	 ("00000000000000000000000000000000"),	 -- 582	0
	 ("00000000000000000000000000000000"),	 -- 581	0
	 ("00000000000000000000000000000000"),	 -- 580	0
	 ("00000000000000000000000000000000"),	 -- 579	0
	 ("00000000000000000000000000000000"),	 -- 578	0
	 ("00000000000000000000000000000000"),	 -- 577	0
	 ("00000000000000000000000000000000"),	 -- 576	0
	 ("00000000000000000000000000000000"),	 -- 575	0
	 ("00000000000000000000000000000000"),	 -- 574	0
	 ("00000000000000000000000000000000"),	 -- 573	0
	 ("00000000000000000000000000000000"),	 -- 572	0
	 ("00000000000000000000000000000000"),	 -- 571	0
	 ("00000000000000000000000000000000"),	 -- 570	0
	 ("00000000000000000000000000000000"),	 -- 569	0
	 ("00000000000000000000000000000000"),	 -- 568	0
	 ("00000000000000000000000000000000"),	 -- 567	0
	 ("00000000000000000000000000000000"),	 -- 566	0
	 ("00000000000000000000000000000000"),	 -- 565	0
	 ("00000000000000000000000000000000"),	 -- 564	0
	 ("00000000000000000000000000000000"),	 -- 563	0
	 ("00000000000000000000000000000000"),	 -- 562	0
	 ("00000000000000000000000000000000"),	 -- 561	0
	 ("00000000000000000000000000000000"),	 -- 560	0
	 ("00000000000000000000000000000000"),	 -- 559	0
	 ("00000000000000000000000000000000"),	 -- 558	0
	 ("00000000000000000000000000000000"),	 -- 557	0
	 ("00000000000000000000000000000000"),	 -- 556	0
	 ("00000000000000000000000000000000"),	 -- 555	0
	 ("00000000000000000000000000000000"),	 -- 554	0
	 ("00000000000000000000000000000000"),	 -- 553	0
	 ("00000000000000000000000000000000"),	 -- 552	0
	 ("00000000000000000000000000000000"),	 -- 551	0
	 ("00000000000000000000000000000000"),	 -- 550	0
	 ("00000000000000000000000000000000"),	 -- 549	0
	 ("00000000000000000000000000000000"),	 -- 548	0
	 ("00000000000000000000000000000000"),	 -- 547	0
	 ("00000000000000000000000000000000"),	 -- 546	0
	 ("00000000000000000000000000000000"),	 -- 545	0
	 ("00000000000000000000000000000000"),	 -- 544	0
	 ("00000000000000000000000000000000"),	 -- 543	0
	 ("00000000000000000000000000000000"),	 -- 542	0
	 ("00000000000000000000000000000000"),	 -- 541	0
	 ("00000000000000000000000000000000"),	 -- 540	0
	 ("00000000000000000000000000000000"),	 -- 539	0
	 ("00000000000000000000000000000000"),	 -- 538	0
	 ("00000000000000000000000000000000"),	 -- 537	0
	 ("00000000000000000000000000000000"),	 -- 536	0
	 ("00000000000000000000000000000000"),	 -- 535	0
	 ("00000000000000000000000000000000"),	 -- 534	0
	 ("00000000000000000000000000000000"),	 -- 533	0
	 ("00000000000000000000000000000000"),	 -- 532	0
	 ("00000000000000000000000000000000"),	 -- 531	0
	 ("00000000000000000000000000000000"),	 -- 530	0
	 ("00000000000000000000000000000000"),	 -- 529	0
	 ("00000000000000000000000000000000"),	 -- 528	0
	 ("00000000000000000000000000000000"),	 -- 527	0
	 ("00000000000000000000000000000000"),	 -- 526	0
	 ("00000000000000000000000000000000"),	 -- 525	0
	 ("00000000000000000000000000000000"),	 -- 524	0
	 ("00000000000000000000000000000000"),	 -- 523	0
	 ("00000000000000000000000000000000"),	 -- 522	0
	 ("00000000000000000000000000000000"),	 -- 521	0
	 ("00000000000000000000000000000000"),	 -- 520	0
	 ("00000000000000000000000000000000"),	 -- 519	0
	 ("00000000000000000000000000000000"),	 -- 518	0
	 ("00000000000000000000000000000000"),	 -- 517	0
	 ("00000000000000000000000000000000"),	 -- 516	0
	 ("00000000000000000000000000000000"),	 -- 515	0
	 ("00000000000000000000000000000000"),	 -- 514	0
	 ("00000000000000000000000000000000"),	 -- 513	0
	 ("00000000000000000000000000000000"),	 -- 512	0
	 ("00000000000000000000000000000000"),	 -- 511	0
	 ("00000000000000000000000000000000"),	 -- 510	0
	 ("00000000000000000000000000000000"),	 -- 509	0
	 ("00000000000000000000000000000000"),	 -- 508	0
	 ("00000000000000000000000000000000"),	 -- 507	0
	 ("00000000000000000000000000000000"),	 -- 506	0
	 ("00000000000000000000000000000000"),	 -- 505	0
	 ("00000000000000000000000000000000"),	 -- 504	0
	 ("00000000000000000000000000000000"),	 -- 503	0
	 ("00000000000000000000000000000000"),	 -- 502	0
	 ("00000000000000000000000000000000"),	 -- 501	0
	 ("00000000000000000000000000000000"),	 -- 500	0
	 ("00000000000000000000000000000000"),	 -- 499	0
	 ("00000000000000000000000000000000"),	 -- 498	0
	 ("00000000000000000000000000000000"),	 -- 497	0
	 ("00000000000000000000000000000000"),	 -- 496	0
	 ("00000000000000000000000000000000"),	 -- 495	0
	 ("00000000000000000000000000000000"),	 -- 494	0
	 ("00000000000000000000000000000000"),	 -- 493	0
	 ("00000000000000000000000000000000"),	 -- 492	0
	 ("00000000000000000000000000000000"),	 -- 491	0
	 ("00000000000000000000000000000000"),	 -- 490	0
	 ("00000000000000000000000000000000"),	 -- 489	0
	 ("00000000000000000000000000000000"),	 -- 488	0
	 ("00000000000000000000000000000000"),	 -- 487	0
	 ("00000000000000000000000000000000"),	 -- 486	0
	 ("00000000000000000000000000000000"),	 -- 485	0
	 ("00000000000000000000000000000000"),	 -- 484	0
	 ("00000000000000000000000000000000"),	 -- 483	0
	 ("00000000000000000000000000000000"),	 -- 482	0
	 ("00000000000000000000000000000000"),	 -- 481	0
	 ("00000000000000000000000000000000"),	 -- 480	0
	 ("00000000000000000000000000000000"),	 -- 479	0
	 ("00000000000000000000000000000000"),	 -- 478	0
	 ("00000000000000000000000000000000"),	 -- 477	0
	 ("00000000000000000000000000000000"),	 -- 476	0
	 ("00000000000000000000000000000000"),	 -- 475	0
	 ("00000000000000000000000000000000"),	 -- 474	0
	 ("00000000000000000000000000000000"),	 -- 473	0
	 ("00000000000000000000000000000000"),	 -- 472	0
	 ("00000000000000000000000000000000"),	 -- 471	0
	 ("00000000000000000000000000000000"),	 -- 470	0
	 ("00000000000000000000000000000000"),	 -- 469	0
	 ("00000000000000000000000000000000"),	 -- 468	0
	 ("00000000000000000000000000000000"),	 -- 467	0
	 ("00000000000000000000000000000000"),	 -- 466	0
	 ("00000000000000000000000000000000"),	 -- 465	0
	 ("00000000000000000000000000000000"),	 -- 464	0
	 ("00000000000000000000000000000000"),	 -- 463	0
	 ("00000000000000000000000000000000"),	 -- 462	0
	 ("00000000000000000000000000000000"),	 -- 461	0
	 ("00000000000000000000000000000000"),	 -- 460	0
	 ("00000000000000000000000000000000"),	 -- 459	0
	 ("00000000000000000000000000000000"),	 -- 458	0
	 ("00000000000000000000000000000000"),	 -- 457	0
	 ("00000000000000000000000000000000"),	 -- 456	0
	 ("00000000000000000000000000000000"),	 -- 455	0
	 ("00000000000000000000000000000000"),	 -- 454	0
	 ("00000000000000000000000000000000"),	 -- 453	0
	 ("00000000000000000000000000000000"),	 -- 452	0
	 ("00000000000000000000000000000000"),	 -- 451	0
	 ("00000000000000000000000000000000"),	 -- 450	0
	 ("00000000000000000000000000000000"),	 -- 449	0
	 ("00000000000000000000000000000000"),	 -- 448	0
	 ("00000000000000000000000000000000"),	 -- 447	0
	 ("00000000000000000000000000000000"),	 -- 446	0
	 ("00000000000000000000000000000000"),	 -- 445	0
	 ("00000000000000000000000000000000"),	 -- 444	0
	 ("00000000000000000000000000000000"),	 -- 443	0
	 ("00000000000000000000000000000000"),	 -- 442	0
	 ("00000000000000000000000000000000"),	 -- 441	0
	 ("00000000000000000000000000000000"),	 -- 440	0
	 ("00000000000000000000000000000000"),	 -- 439	0
	 ("00000000000000000000000000000000"),	 -- 438	0
	 ("00000000000000000000000000000000"),	 -- 437	0
	 ("00000000000000000000000000000000"),	 -- 436	0
	 ("00000000000000000000000000000000"),	 -- 435	0
	 ("00000000000000000000000000000000"),	 -- 434	0
	 ("00000000000000000000000000000000"),	 -- 433	0
	 ("00000000000000000000000000000000"),	 -- 432	0
	 ("00000000000000000000000000000000"),	 -- 431	0
	 ("00000000000000000000000000000000"),	 -- 430	0
	 ("00000000000000000000000000000000"),	 -- 429	0
	 ("00000000000000000000000000000000"),	 -- 428	0
	 ("00000000000000000000000000000000"),	 -- 427	0
	 ("00000000000000000000000000000000"),	 -- 426	0
	 ("00000000000000000000000000000000"),	 -- 425	0
	 ("00000000000000000000000000000000"),	 -- 424	0
	 ("00000000000000000000000000000000"),	 -- 423	0
	 ("00000000000000000000000000000000"),	 -- 422	0
	 ("00000000000000000000000000000000"),	 -- 421	0
	 ("00000000000000000000000000000000"),	 -- 420	0
	 ("00000000000000000000000000000000"),	 -- 419	0
	 ("00000000000000000000000000000000"),	 -- 418	0
	 ("00000000000000000000000000000000"),	 -- 417	0
	 ("00000000000000000000000000000000"),	 -- 416	0
	 ("00000000000000000000000000000000"),	 -- 415	0
	 ("00000000000000000000000000000000"),	 -- 414	0
	 ("00000000000000000000000000000000"),	 -- 413	0
	 ("00000000000000000000000000000000"),	 -- 412	0
	 ("00000000000000000000000000000000"),	 -- 411	0
	 ("00000000000000000000000000000000"),	 -- 410	0
	 ("00000000000000000000000000000000"),	 -- 409	0
	 ("00000000000000000000000000000000"),	 -- 408	0
	 ("00000000000000000000000000000000"),	 -- 407	0
	 ("00000000000000000000000000000000"),	 -- 406	0
	 ("00000000000000000000000000000000"),	 -- 405	0
	 ("00000000000000000000000000000000"),	 -- 404	0
	 ("00000000000000000000000000000000"),	 -- 403	0
	 ("00000000000000000000000000000000"),	 -- 402	0
	 ("00000000000000000000000000000000"),	 -- 401	0
	 ("00000000000000000000000000000000"),	 -- 400	0
	 ("00000000000000000000000000000000"),	 -- 399	0
	 ("00000000000000000000000000000000"),	 -- 398	0
	 ("00000000000000000000000000000000"),	 -- 397	0
	 ("00000000000000000000000000000000"),	 -- 396	0
	 ("00000000000000000000000000000000"),	 -- 395	0
	 ("00000000000000000000000000000000"),	 -- 394	0
	 ("00000000000000000000000000000000"),	 -- 393	0
	 ("00000000000000000000000000000000"),	 -- 392	0
	 ("00000000000000000000000000000000"),	 -- 391	0
	 ("00000000000000000000000000000000"),	 -- 390	0
	 ("00000000000000000000000000000000"),	 -- 389	0
	 ("00000000000000000000000000000000"),	 -- 388	0
	 ("00000000000000000000000000000000"),	 -- 387	0
	 ("00000000000000000000000000000000"),	 -- 386	0
	 ("00000000000000000000000000000000"),	 -- 385	0
	 ("00000000000000000000000000000000"),	 -- 384	0
	 ("00000000000000000000000000000000"),	 -- 383	0
	 ("00000000000000000000000000000000"),	 -- 382	0
	 ("00000000000000000000000000000000"),	 -- 381	0
	 ("00000000000000000000000000000000"),	 -- 380	0
	 ("00000000000000000000000000000000"),	 -- 379	0
	 ("00000000000000000000000000000000"),	 -- 378	0
	 ("00000000000000000000000000000000"),	 -- 377	0
	 ("00000000000000000000000000000000"),	 -- 376	0
	 ("00000000000000000000000000000000"),	 -- 375	0
	 ("00000000000000000000000000000000"),	 -- 374	0
	 ("00000000000000000000000000000000"),	 -- 373	0
	 ("00000000000000000000000000000000"),	 -- 372	0
	 ("00000000000000000000000000000000"),	 -- 371	0
	 ("00000000000000000000000000000000"),	 -- 370	0
	 ("00000000000000000000000000000000"),	 -- 369	0
	 ("00000000000000000000000000000000"),	 -- 368	0
	 ("00000000000000000000000000000000"),	 -- 367	0
	 ("00000000000000000000000000000000"),	 -- 366	0
	 ("00000000000000000000000000000000"),	 -- 365	0
	 ("00000000000000000000000000000000"),	 -- 364	0
	 ("00000000000000000000000000000000"),	 -- 363	0
	 ("00000000000000000000000000000000"),	 -- 362	0
	 ("00000000000000000000000000000000"),	 -- 361	0
	 ("00000000000000000000000000000000"),	 -- 360	0
	 ("00000000000000000000000000000000"),	 -- 359	0
	 ("00000000000000000000000000000000"),	 -- 358	0
	 ("00000000000000000000000000000000"),	 -- 357	0
	 ("00000000000000000000000000000000"),	 -- 356	0
	 ("00000000000000000000000000000000"),	 -- 355	0
	 ("00000000000000000000000000000000"),	 -- 354	0
	 ("00000000000000000000000000000000"),	 -- 353	0
	 ("00000000000000000000000000000000"),	 -- 352	0
	 ("00000000000000000000000000000000"),	 -- 351	0
	 ("00000000000000000000000000000000"),	 -- 350	0
	 ("00000000000000000000000000000000"),	 -- 349	0
	 ("00000000000000000000000000000000"),	 -- 348	0
	 ("00000000000000000000000000000000"),	 -- 347	0
	 ("00000000000000000000000000000000"),	 -- 346	0
	 ("00000000000000000000000000000000"),	 -- 345	0
	 ("00000000000000000000000000000000"),	 -- 344	0
	 ("00000000000000000000000000000000"),	 -- 343	0
	 ("00000000000000000000000000000000"),	 -- 342	0
	 ("00000000000000000000000000000000"),	 -- 341	0
	 ("00000000000000000000000000000000"),	 -- 340	0
	 ("00000000000000000000000000000000"),	 -- 339	0
	 ("00000000000000000000000000000000"),	 -- 338	0
	 ("00000000000000000000000000000000"),	 -- 337	0
	 ("00000000000000000000000000000000"),	 -- 336	0
	 ("00000000000000000000000000000000"),	 -- 335	0
	 ("00000000000000000000000000000000"),	 -- 334	0
	 ("00000000000000000000000000000000"),	 -- 333	0
	 ("00000000000000000000000000000000"),	 -- 332	0
	 ("00000000000000000000000000000000"),	 -- 331	0
	 ("00000000000000000000000000000000"),	 -- 330	0
	 ("00000000000000000000000000000000"),	 -- 329	0
	 ("00000000000000000000000000000000"),	 -- 328	0
	 ("00000000000000000000000000000000"),	 -- 327	0
	 ("00000000000000000000000000000000"),	 -- 326	0
	 ("00000000000000000000000000000000"),	 -- 325	0
	 ("00000000000000000000000000000000"),	 -- 324	0
	 ("00000000000000000000000000000000"),	 -- 323	0
	 ("00000000000000000000000000000000"),	 -- 322	0
	 ("00000000000000000000000000000000"),	 -- 321	0
	 ("00000000000000000000000000000000"),	 -- 320	0
	 ("00000000000000000000000000000000"),	 -- 319	0
	 ("00000000000000000000000000000000"),	 -- 318	0
	 ("00000000000000000000000000000000"),	 -- 317	0
	 ("00000000000000000000000000000000"),	 -- 316	0
	 ("00000000000000000000000000000000"),	 -- 315	0
	 ("00000000000000000000000000000000"),	 -- 314	0
	 ("00000000000000000000000000000000"),	 -- 313	0
	 ("00000000000000000000000000000000"),	 -- 312	0
	 ("00000000000000000000000000000000"),	 -- 311	0
	 ("00000000000000000000000000000000"),	 -- 310	0
	 ("00000000000000000000000000000000"),	 -- 309	0
	 ("00000000000000000000000000000000"),	 -- 308	0
	 ("00000000000000000000000000000000"),	 -- 307	0
	 ("00000000000000000000000000000000"),	 -- 306	0
	 ("00000000000000000000000000000000"),	 -- 305	0
	 ("00000000000000000000000000000000"),	 -- 304	0
	 ("00000000000000000000000000000000"),	 -- 303	0
	 ("00000000000000000000000000000000"),	 -- 302	0
	 ("00000000000000000000000000000000"),	 -- 301	0
	 ("00000000000000000000000000000000"),	 -- 300	0
	 ("00000000000000000000000000000000"),	 -- 299	0
	 ("00000000000000000000000000000000"),	 -- 298	0
	 ("00000000000000000000000000000000"),	 -- 297	0
	 ("00000000000000000000000000000000"),	 -- 296	0
	 ("00000000000000000000000000000000"),	 -- 295	0
	 ("00000000000000000000000000000000"),	 -- 294	0
	 ("00000000000000000000000000000000"),	 -- 293	0
	 ("00000000000000000000000000000000"),	 -- 292	0
	 ("00000000000000000000000000000000"),	 -- 291	0
	 ("00000000000000000000000000000000"),	 -- 290	0
	 ("00000000000000000000000000000000"),	 -- 289	0
	 ("00000000000000000000000000000000"),	 -- 288	0
	 ("00000000000000000000000000000000"),	 -- 287	0
	 ("00000000000000000000000000000000"),	 -- 286	0
	 ("00000000000000000000000000000000"),	 -- 285	0
	 ("00000000000000000000000000000000"),	 -- 284	0
	 ("00000000000000000000000000000000"),	 -- 283	0
	 ("00000000000000000000000000000000"),	 -- 282	0
	 ("00000000000000000000000000000000"),	 -- 281	0
	 ("00000000000000000000000000000000"),	 -- 280	0
	 ("00000000000000000000000000000000"),	 -- 279	0
	 ("00000000000000000000000000000000"),	 -- 278	0
	 ("00000000000000000000000000000000"),	 -- 277	0
	 ("00000000000000000000000000000000"),	 -- 276	0
	 ("00000000000000000000000000000000"),	 -- 275	0
	 ("00000000000000000000000000000000"),	 -- 274	0
	 ("00000000000000000000000000000000"),	 -- 273	0
	 ("00000000000000000000000000000000"),	 -- 272	0
	 ("00000000000000000000000000000000"),	 -- 271	0
	 ("00000000000000000000000000000000"),	 -- 270	0
	 ("00000000000000000000000000000000"),	 -- 269	0
	 ("00000000000000000000000000000000"),	 -- 268	0
	 ("00000000000000000000000000000000"),	 -- 267	0
	 ("00000000000000000000000000000000"),	 -- 266	0
	 ("00000000000000000000000000000000"),	 -- 265	0
	 ("00000000000000000000000000000000"),	 -- 264	0
	 ("00000000000000000000000000000000"),	 -- 263	0
	 ("00000000000000000000000000000000"),	 -- 262	0
	 ("00000000000000000000000000000000"),	 -- 261	0
	 ("00000000000000000000000000000000"),	 -- 260	0
	 ("00000000000000000000000000000000"),	 -- 259	0
	 ("00000000000000000000000000000000"),	 -- 258	0
	 ("00000000000000000000000000000000"),	 -- 257	0
	 ("00000000000000000000000000000000"),	 -- 256	0
	 ("00000000000000000000000000000000"),	 -- 255	0
	 ("00000000000000000000000000000000"),	 -- 254	0
	 ("00000000000000000000000000000000"),	 -- 253	0
	 ("00000000000000000000000000000000"),	 -- 252	0
	 ("00000000000000000000000000000000"),	 -- 251	0
	 ("00000000000000000000000000000000"),	 -- 250	0
	 ("00000000000000000000000000000000"),	 -- 249	0
	 ("00000000000000000000000000000000"),	 -- 248	0
	 ("00000000000000000000000000000000"),	 -- 247	0
	 ("00000000000000000000000000000000"),	 -- 246	0
	 ("00000000000000000000000000000000"),	 -- 245	0
	 ("00000000000000000000000000000000"),	 -- 244	0
	 ("00000000000000000000000000000000"),	 -- 243	0
	 ("00000000000000000000000000000000"),	 -- 242	0
	 ("00000000000000000000000000000000"),	 -- 241	0
	 ("00000000000000000000000000000000"),	 -- 240	0
	 ("00000000000000000000000000000000"),	 -- 239	0
	 ("00000000000000000000000000000000"),	 -- 238	0
	 ("00000000000000000000000000000000"),	 -- 237	0
	 ("00000000000000000000000000000000"),	 -- 236	0
	 ("00000000000000000000000000000000"),	 -- 235	0
	 ("00000000000000000000000000000000"),	 -- 234	0
	 ("00000000000000000000000000000000"),	 -- 233	0
	 ("00000000000000000000000000000000"),	 -- 232	0
	 ("00000000000000000000000000000000"),	 -- 231	0
	 ("00000000000000000000000000000000"),	 -- 230	0
	 ("00000000000000000000000000000000"),	 -- 229	0
	 ("00000000000000000000000000000000"),	 -- 228	0
	 ("00000000000000000000000000000000"),	 -- 227	0
	 ("00000000000000000000000000000000"),	 -- 226	0
	 ("00000000000000000000000000000000"),	 -- 225	0
	 ("00000000000000000000000000000000"),	 -- 224	0
	 ("00000000000000000000000000000000"),	 -- 223	0
	 ("00000000000000000000000000000000"),	 -- 222	0
	 ("00000000000000000000000000000000"),	 -- 221	0
	 ("00000000000000000000000000000000"),	 -- 220	0
	 ("00000000000000000000000000000000"),	 -- 219	0
	 ("00000000000000000000000000000000"),	 -- 218	0
	 ("00000000000000000000000000000000"),	 -- 217	0
	 ("00000000000000000000000000000000"),	 -- 216	0
	 ("00000000000000000000000000000000"),	 -- 215	0
	 ("00000000000000000000000000000000"),	 -- 214	0
	 ("00000000000000000000000000000000"),	 -- 213	0
	 ("00000000000000000000000000000000"),	 -- 212	0
	 ("00000000000000000000000000000000"),	 -- 211	0
	 ("00000000000000000000000000000000"),	 -- 210	0
	 ("00000000000000000000000000000000"),	 -- 209	0
	 ("00000000000000000000000000000000"),	 -- 208	0
	 ("00000000000000000000000000000000"),	 -- 207	0
	 ("00000000000000000000000000000000"),	 -- 206	0
	 ("00000000000000000000000000000000"),	 -- 205	0
	 ("00000000000000000000000000000000"),	 -- 204	0
	 ("00000000000000000000000000000000"),	 -- 203	0
	 ("00000000000000000000000000000000"),	 -- 202	0
	 ("00000000000000000000000000000000"),	 -- 201	0
	 ("00000000000000000000000000000000"),	 -- 200	0
	 ("00000000000000000000000000000000"),	 -- 199	0
	 ("00000000000000000000000000000000"),	 -- 198	0
	 ("00000000000000000000000000000000"),	 -- 197	0
	 ("00000000000000000000000000000000"),	 -- 196	0
	 ("00000000000000000000000000000000"),	 -- 195	0
	 ("00000000000000000000000000000000"),	 -- 194	0
	 ("00000000000000000000000000000000"),	 -- 193	0
	 ("00000000000000000000000000000000"),	 -- 192	0
	 ("00000000000000000000000000000000"),	 -- 191	0
	 ("00000000000000000000000000000000"),	 -- 190	0
	 ("00000000000000000000000000000000"),	 -- 189	0
	 ("00000000000000000000000000000000"),	 -- 188	0
	 ("00000000000000000000000000000000"),	 -- 187	0
	 ("00000000000000000000000000000000"),	 -- 186	0
	 ("00000000000000000000000000000000"),	 -- 185	0
	 ("00000000000000000000000000000000"),	 -- 184	0
	 ("00000000000000000000000000000000"),	 -- 183	0
	 ("00000000000000000000000000000000"),	 -- 182	0
	 ("00000000000000000000000000000000"),	 -- 181	0
	 ("00000000000000000000000000000000"),	 -- 180	0
	 ("00000000000000000000000000000000"),	 -- 179	0
	 ("00000000000000000000000000000000"),	 -- 178	0
	 ("00000000000000000000000000000000"),	 -- 177	0
	 ("00000000000000000000000000000000"),	 -- 176	0
	 ("00000000000000000000000000000000"),	 -- 175	0
	 ("00000000000000000000000000000000"),	 -- 174	0
	 ("00000000000000000000000000000000"),	 -- 173	0
	 ("00000000000000000000000000000000"),	 -- 172	0
	 ("00000000000000000000000000000000"),	 -- 171	0
	 ("00000000000000000000000000000000"),	 -- 170	0
	 ("00000000000000000000000000000000"),	 -- 169	0
	 ("00000000000000000000000000000000"),	 -- 168	0
	 ("00000000000000000000000000000000"),	 -- 167	0
	 ("00000000000000000000000000000000"),	 -- 166	0
	 ("00000000000000000000000000000000"),	 -- 165	0
	 ("00000000000000000000000000000000"),	 -- 164	0
	 ("00000000000000000000000000000000"),	 -- 163	0
	 ("00000000000000000000000000000000"),	 -- 162	0
	 ("00000000000000000000000000000000"),	 -- 161	0
	 ("00000000000000000000000000000000"),	 -- 160	0
	 ("00000000000000000000000000000000"),	 -- 159	0
	 ("00000000000000000000000000000000"),	 -- 158	0
	 ("00000000000000000000000000000000"),	 -- 157	0
	 ("00000000000000000000000000000000"),	 -- 156	0
	 ("00000000000000000000000000000000"),	 -- 155	0
	 ("00000000000000000000000000000000"),	 -- 154	0
	 ("00000000000000000000000000000000"),	 -- 153	0
	 ("00000000000000000000000000000000"),	 -- 152	0
	 ("00000000000000000000000000000000"),	 -- 151	0
	 ("00000000000000000000000000000000"),	 -- 150	0
	 ("00000000000000000000000000000000"),	 -- 149	0
	 ("00000000000000000000000000000000"),	 -- 148	0
	 ("00000000000000000000000000000000"),	 -- 147	0
	 ("00000000000000000000000000000000"),	 -- 146	0
	 ("00000000000000000000000000000000"),	 -- 145	0
	 ("00000000000000000000000000000000"),	 -- 144	0
	 ("00000000000000000000000000000000"),	 -- 143	0
	 ("00000000000000000000000000000000"),	 -- 142	0
	 ("00000000000000000000000000000000"),	 -- 141	0
	 ("00000000000000000000000000000000"),	 -- 140	0
	 ("00000000000000000000000000000000"),	 -- 139	0
	 ("00000000000000000000000000000000"),	 -- 138	0
	 ("00000000000000000000000000000000"),	 -- 137	0
	 ("00000000000000000000000000000000"),	 -- 136	0
	 ("00000000000000000000000000000000"),	 -- 135	0
	 ("00000000000000000000000000000000"),	 -- 134	0
	 ("00000000000000000000000000000000"),	 -- 133	0
	 ("00000000000000000000000000000000"),	 -- 132	0
	 ("00000000000000000000000000000000"),	 -- 131	0
	 ("00000000000000000000000000000000"),	 -- 130	0
	 ("00000000000000000000000000000000"),	 -- 129	0
	 ("00000000000000000000000000000000"),	 -- 128	0
	 ("00000000000000000000000000000000"),	 -- 127	0
	 ("00000000000000000000000000000000"),	 -- 126	0
	 ("00000000000000000000000000000000"),	 -- 125	0
	 ("00000000000000000000000000000000"),	 -- 124	0
	 ("00000000000000000000000000000000"),	 -- 123	0
	 ("00000000000000000000000000000000"),	 -- 122	0
	 ("00000000000000000000000000000000"),	 -- 121	0
	 ("00000000000000000000000000000000"),	 -- 120	0
	 ("00000000000000000000000000000000"),	 -- 119	0
	 ("00000000000000000000000000000000"),	 -- 118	0
	 ("00000000000000000000000000000000"),	 -- 117	0
	 ("00000000000000000000000000000000"),	 -- 116	0
	 ("00000000000000000000000000000000"),	 -- 115	0
	 ("00000000000000000000000000000000"),	 -- 114	0
	 ("00000000000000000000000000000000"),	 -- 113	0
	 ("00000000000000000000000000000000"),	 -- 112	0
	 ("00000000000000000000000000000000"),	 -- 111	0
	 ("00000000000000000000000000000000"),	 -- 110	0
	 ("00000000000000000000000000000000"),	 -- 109	0
	 ("00000000000000000000000000000000"),	 -- 108	0
	 ("00000000000000000000000000000000"),	 -- 107	0
	 ("00000000000000000000000000000000"),	 -- 106	0
	 ("00000000000000000000000000000000"),	 -- 105	0
	 ("00000000000000000000000000000000"),	 -- 104	0
	 ("00000000000000000000000000000000"),	 -- 103	0
	 ("00000000000000000000000000000000"),	 -- 102	0
	 ("00000000000000000000000000000000"),	 -- 101	0
	 ("00000000000000000000000000000000"),	 -- 100	0
	 ("00000000000000000000000000000000"),	 -- 99	0
	 ("00000000000000000000000000000000"),	 -- 98	0
	 ("00000000000000000000000000000000"),	 -- 97	0
	 ("00000000000000000000000000000000"),	 -- 96	0
	 ("00000000000000000000000000000000"),	 -- 95	0
	 ("00000000000000000000000000000000"),	 -- 94	0
	 ("00000000000000000000000000000000"),	 -- 93	0
	 ("00000000000000000000000000000000"),	 -- 92	0
	 ("00000000000000000000000000000000"),	 -- 91	0
	 ("00000000000000000000000000000000"),	 -- 90	0
	 ("00000000000000000000000000000000"),	 -- 89	0
	 ("00000000000000000000000000000000"),	 -- 88	0
	 ("00000000000000000000000000000000"),	 -- 87	0
	 ("00000000000000000000000000000000"),	 -- 86	0
	 ("00000000000000000000000000000000"),	 -- 85	0
	 ("00000000000000000000000000000000"),	 -- 84	0
	 ("00000000000000000000000000000000"),	 -- 83	0
	 ("00000000000000000000000000000000"),	 -- 82	0
	 ("00000000000000000000000000000000"),	 -- 81	0
	 ("00000000000000000000000000000000"),	 -- 80	0
	 ("00000000000000000000000000000000"),	 -- 79	0
	 ("00000000000000000000000000000000"),	 -- 78	0
	 ("00000000000000000000000000000000"),	 -- 77	0
	 ("00000000000000000000000000000000"),	 -- 76	0
	 ("00000000000000000000000000000000"),	 -- 75	0
	 ("00000000000000000000000000000000"),	 -- 74	0
	 ("00000000000000000000000000000000"),	 -- 73	0
	 ("00000000000000000000000000000000"),	 -- 72	0
	 ("00000000000000000000000000000000"),	 -- 71	0
	 ("00000000000000000000000000000000"),	 -- 70	0
	 ("00000000000000000000000000000000"),	 -- 69	0
	 ("00000000000000000000000000000000"),	 -- 68	0
	 ("00000000000000000000000000000000"),	 -- 67	0
	 ("00000000000000000000000000000000"),	 -- 66	0
	 ("00000000000000000000000000000000"),	 -- 65	0
	 ("00000000000000000000000000000000"),	 -- 64	0
	 ("00000000000000000000000000000000"),	 -- 63	0
	 ("00000000000000000000000000000000"),	 -- 62	0
	 ("00000000000000000000000000000000"),	 -- 61	0
	 ("00000000000000000000000000000000"),	 -- 60	0
	 ("00000000000000000000000000000000"),	 -- 59	0
	 ("00000000000000000000000000000000"),	 -- 58	0
	 ("00000000000000000000000000000000"),	 -- 57	0
	 ("00000000000000000000000000000000"),	 -- 56	0
	 ("00000000000000000000000000000000"),	 -- 55	0
	 ("00000000000000000000000000000000"),	 -- 54	0
	 ("00000000000000000000000000000000"),	 -- 53	0
	 ("00000000000000000000000000000000"),	 -- 52	0
	 ("00000000000000000000000000000000"),	 -- 51	0
	 ("00000000000000000000000000000000"),	 -- 50	0
	 ("00000000000000000000000000000000"),	 -- 49	0
	 ("00000000000000000000000000000000"),	 -- 48	0
	 ("00000000000000000000000000000000"),	 -- 47	0
	 ("00000000000000000000000000000000"),	 -- 46	0
	 ("00000000000000000000000000000000"),	 -- 45	0
	 ("00000000000000000000000000000000"),	 -- 44	0
	 ("00000000000000000000000000000000"),	 -- 43	0
	 ("00000000000000000000000000000000"),	 -- 42	0
	 ("00000000000000000000000000000000"),	 -- 41	0
	 ("00000000000000000000000000000000"),	 -- 40	0
	 ("00000000000000000000000000000000"),	 -- 39	0
	 ("00000000000000000000000000000000"),	 -- 38	0
	 ("00000000000000000000000000000000"),	 -- 37	0
	 ("00000000000000000000000000000000"),	 -- 36	0
	 ("00000000000000000000000000000000"),	 -- 35	0
	 ("00000000000000000000000000000000"),	 -- 34	0
	 ("00000000000000000000000000000000"),	 -- 33	0
	 ("00000000000000000000000000000000"),	 -- 32	0
	 ("00000000000000000000000000000000"),	 -- 31	0
	 ("00000000000000000000000000000000"),	 -- 30	0
	 ("00000000000000000000000000000000"),	 -- 29	0
	 ("00000000000000000000000000000000"),	 -- 28	0
	 ("00000000000000000000000000000000"),	 -- 27	0
	 ("00000000000000000000000000000000"),	 -- 26	0
	 ("00000000000000000000000000000000"),	 -- 25	0
	 ("00000000000000000000000000000000"),	 -- 24	0
	 ("00000000000000000000000000000000"),	 -- 23	0
	 ("00000000000000000000000000000000"),	 -- 22	0
	 ("00000000000000000000000000000000"),	 -- 21	0
	 ("00000000000000000000000000000000"),	 -- 20	0
	 ("00000000000000000000000000000000"),	 -- 19	0
	 ("00000000000000000000000000000000"),	 -- 18	0
	 ("00000000000000000000000000000000"),	 -- 17	0
	 ("00000000000000000000000000000000"),	 -- 16	0
	 ("00000000000000000000000000000000"),	 -- 15	0
	 ("00000000000000000000000000000000"),	 -- 14	0
	 ("00000000000000000000000000000000"),	 -- 13	0
	 ("00000000000000000000000000000000"),	 -- 12	0
	 ("00000000000000000000000000000000"),	 -- 11	0
	 ("00000000000000000000000000000000"),	 -- 10	0
	 ("00000000000000000000000000000000"),	 -- 9	0
	 ("00000000000000000000000000000000"),	 -- 8	0
	 ("00000000000000000000000000000000"),	 -- 7	0
	 ("00000000000000000000000000000000"),	 -- 6	0
	 ("00000000000000000000000000000000"),	 -- 5	0
	 ("00000000000000000000000000000000"),	 -- 4	0
	 ("00000000000000000000000000000000"),	 -- 3	0
	 ("00000000000000000000000000000011"),	 -- 2	3
	 ("00000000000000000000000000000010"),	 -- 1	2
	 ("00000000000000000000000000000001"));	 -- 0	1


begin 
       process (clk) 
       begin 
              if (clk'event and clk = '1') then 
                  if (we_0 = '1') then 
                        RAM(conv_integer(address_0)) <= data_in_0; 
                        data_out_0 <= RAM(conv_integer(read_a)); 
                  elsif (oe_0 = '1') then 
                        data_out_0 <= RAM(conv_integer(read_a)); 
                  end if; 
                  read_a <= address_0; 
             end if; 
       end process; 
       process (clk) 
       begin 
              if (clk'event and clk = '1') then 
                  if (we_1 = '1') then 
                        RAM(conv_integer(address_1)) <= data_in_1; 
                        data_out_1 <= RAM(conv_integer(read_b)); 
                  elsif (oe_1 = '1') then 
                        data_out_1 <= RAM(conv_integer(read_b)); 
                  end if; 
                  read_b <= address_1; 
             end if; 
       end process; 
end rtl; 

library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 

entity dual_block_ram_y is 
generic( 
	data_width : integer := 8; 
	address_width : integer := 8 
); 
port( 
	data_in_0 : in std_logic_vector(data_width-1 downto 0) := (others => '0'); 
	address_0 : in std_logic_vector(address_width-1 downto 0); 
	we_0: in std_logic := '0'; 
	oe_0: in std_logic := '1'; 
	data_out_0 : out std_logic_vector(data_width-1 downto 0); 
	data_in_1 : in std_logic_vector(data_width-1 downto 0) := (others => '0'); 
	address_1 : in std_logic_vector(address_width-1 downto 0); 
	we_1: in std_logic := '0'; 
	oe_1: in std_logic := '1'; 
	data_out_1 : out std_logic_vector(data_width-1 downto 0); 
	clk : in std_logic); 
end dual_block_ram_y; 

architecture rtl of dual_block_ram_y is 

constant mem_depth : integer := 2**address_width; 
type ram_type is array (mem_depth-1 downto 0) 
of std_logic_vector (data_width-1 downto 0); 

signal read_a : std_logic_vector(address_width-1 downto 0); 
signal read_b : std_logic_vector(address_width-1 downto 0); 
signal RAM : ram_type := ram_type'( 
	 ("00000000000000000000000000000101"),	 -- 2047	5
	 ("00000000000000000000000000000000"),	 -- 2046	0
	 ("00000000000000000000000000000000"),	 -- 2045	0
	 ("00000000000000000000000000000000"),	 -- 2044	0
	 ("00000000000000000000000000000000"),	 -- 2043	0
	 ("00000000000000000000000000000000"),	 -- 2042	0
	 ("00000000000000000000000000000000"),	 -- 2041	0
	 ("00000000000000000000000000000000"),	 -- 2040	0
	 ("00000000000000000000000000000000"),	 -- 2039	0
	 ("00000000000000000000000000000000"),	 -- 2038	0
	 ("00000000000000000000000000000000"),	 -- 2037	0
	 ("00000000000000000000000000000000"),	 -- 2036	0
	 ("00000000000000000000000000000000"),	 -- 2035	0
	 ("00000000000000000000000000000000"),	 -- 2034	0
	 ("00000000000000000000000000000000"),	 -- 2033	0
	 ("00000000000000000000000000000000"),	 -- 2032	0
	 ("00000000000000000000000000000000"),	 -- 2031	0
	 ("00000000000000000000000000000000"),	 -- 2030	0
	 ("00000000000000000000000000000000"),	 -- 2029	0
	 ("00000000000000000000000000000000"),	 -- 2028	0
	 ("00000000000000000000000000000000"),	 -- 2027	0
	 ("00000000000000000000000000000000"),	 -- 2026	0
	 ("00000000000000000000000000000000"),	 -- 2025	0
	 ("00000000000000000000000000000000"),	 -- 2024	0
	 ("00000000000000000000000000000000"),	 -- 2023	0
	 ("00000000000000000000000000000000"),	 -- 2022	0
	 ("00000000000000000000000000000000"),	 -- 2021	0
	 ("00000000000000000000000000000000"),	 -- 2020	0
	 ("00000000000000000000000000000000"),	 -- 2019	0
	 ("00000000000000000000000000000000"),	 -- 2018	0
	 ("00000000000000000000000000000000"),	 -- 2017	0
	 ("00000000000000000000000000000000"),	 -- 2016	0
	 ("00000000000000000000000000000000"),	 -- 2015	0
	 ("00000000000000000000000000000000"),	 -- 2014	0
	 ("00000000000000000000000000000000"),	 -- 2013	0
	 ("00000000000000000000000000000000"),	 -- 2012	0
	 ("00000000000000000000000000000000"),	 -- 2011	0
	 ("00000000000000000000000000000000"),	 -- 2010	0
	 ("00000000000000000000000000000000"),	 -- 2009	0
	 ("00000000000000000000000000000000"),	 -- 2008	0
	 ("00000000000000000000000000000000"),	 -- 2007	0
	 ("00000000000000000000000000000000"),	 -- 2006	0
	 ("00000000000000000000000000000000"),	 -- 2005	0
	 ("00000000000000000000000000000000"),	 -- 2004	0
	 ("00000000000000000000000000000000"),	 -- 2003	0
	 ("00000000000000000000000000000000"),	 -- 2002	0
	 ("00000000000000000000000000000000"),	 -- 2001	0
	 ("00000000000000000000000000000000"),	 -- 2000	0
	 ("00000000000000000000000000000000"),	 -- 1999	0
	 ("00000000000000000000000000000000"),	 -- 1998	0
	 ("00000000000000000000000000000000"),	 -- 1997	0
	 ("00000000000000000000000000000000"),	 -- 1996	0
	 ("00000000000000000000000000000000"),	 -- 1995	0
	 ("00000000000000000000000000000000"),	 -- 1994	0
	 ("00000000000000000000000000000000"),	 -- 1993	0
	 ("00000000000000000000000000000000"),	 -- 1992	0
	 ("00000000000000000000000000000000"),	 -- 1991	0
	 ("00000000000000000000000000000000"),	 -- 1990	0
	 ("00000000000000000000000000000000"),	 -- 1989	0
	 ("00000000000000000000000000000000"),	 -- 1988	0
	 ("00000000000000000000000000000000"),	 -- 1987	0
	 ("00000000000000000000000000000000"),	 -- 1986	0
	 ("00000000000000000000000000000000"),	 -- 1985	0
	 ("00000000000000000000000000000000"),	 -- 1984	0
	 ("00000000000000000000000000000000"),	 -- 1983	0
	 ("00000000000000000000000000000000"),	 -- 1982	0
	 ("00000000000000000000000000000000"),	 -- 1981	0
	 ("00000000000000000000000000000000"),	 -- 1980	0
	 ("00000000000000000000000000000000"),	 -- 1979	0
	 ("00000000000000000000000000000000"),	 -- 1978	0
	 ("00000000000000000000000000000000"),	 -- 1977	0
	 ("00000000000000000000000000000000"),	 -- 1976	0
	 ("00000000000000000000000000000000"),	 -- 1975	0
	 ("00000000000000000000000000000000"),	 -- 1974	0
	 ("00000000000000000000000000000000"),	 -- 1973	0
	 ("00000000000000000000000000000000"),	 -- 1972	0
	 ("00000000000000000000000000000000"),	 -- 1971	0
	 ("00000000000000000000000000000000"),	 -- 1970	0
	 ("00000000000000000000000000000000"),	 -- 1969	0
	 ("00000000000000000000000000000000"),	 -- 1968	0
	 ("00000000000000000000000000000000"),	 -- 1967	0
	 ("00000000000000000000000000000000"),	 -- 1966	0
	 ("00000000000000000000000000000000"),	 -- 1965	0
	 ("00000000000000000000000000000000"),	 -- 1964	0
	 ("00000000000000000000000000000000"),	 -- 1963	0
	 ("00000000000000000000000000000000"),	 -- 1962	0
	 ("00000000000000000000000000000000"),	 -- 1961	0
	 ("00000000000000000000000000000000"),	 -- 1960	0
	 ("00000000000000000000000000000000"),	 -- 1959	0
	 ("00000000000000000000000000000000"),	 -- 1958	0
	 ("00000000000000000000000000000000"),	 -- 1957	0
	 ("00000000000000000000000000000000"),	 -- 1956	0
	 ("00000000000000000000000000000000"),	 -- 1955	0
	 ("00000000000000000000000000000000"),	 -- 1954	0
	 ("00000000000000000000000000000000"),	 -- 1953	0
	 ("00000000000000000000000000000000"),	 -- 1952	0
	 ("00000000000000000000000000000000"),	 -- 1951	0
	 ("00000000000000000000000000000000"),	 -- 1950	0
	 ("00000000000000000000000000000000"),	 -- 1949	0
	 ("00000000000000000000000000000000"),	 -- 1948	0
	 ("00000000000000000000000000000000"),	 -- 1947	0
	 ("00000000000000000000000000000000"),	 -- 1946	0
	 ("00000000000000000000000000000000"),	 -- 1945	0
	 ("00000000000000000000000000000000"),	 -- 1944	0
	 ("00000000000000000000000000000000"),	 -- 1943	0
	 ("00000000000000000000000000000000"),	 -- 1942	0
	 ("00000000000000000000000000000000"),	 -- 1941	0
	 ("00000000000000000000000000000000"),	 -- 1940	0
	 ("00000000000000000000000000000000"),	 -- 1939	0
	 ("00000000000000000000000000000000"),	 -- 1938	0
	 ("00000000000000000000000000000000"),	 -- 1937	0
	 ("00000000000000000000000000000000"),	 -- 1936	0
	 ("00000000000000000000000000000000"),	 -- 1935	0
	 ("00000000000000000000000000000000"),	 -- 1934	0
	 ("00000000000000000000000000000000"),	 -- 1933	0
	 ("00000000000000000000000000000000"),	 -- 1932	0
	 ("00000000000000000000000000000000"),	 -- 1931	0
	 ("00000000000000000000000000000000"),	 -- 1930	0
	 ("00000000000000000000000000000000"),	 -- 1929	0
	 ("00000000000000000000000000000000"),	 -- 1928	0
	 ("00000000000000000000000000000000"),	 -- 1927	0
	 ("00000000000000000000000000000000"),	 -- 1926	0
	 ("00000000000000000000000000000000"),	 -- 1925	0
	 ("00000000000000000000000000000000"),	 -- 1924	0
	 ("00000000000000000000000000000000"),	 -- 1923	0
	 ("00000000000000000000000000000000"),	 -- 1922	0
	 ("00000000000000000000000000000000"),	 -- 1921	0
	 ("00000000000000000000000000000000"),	 -- 1920	0
	 ("00000000000000000000000000000000"),	 -- 1919	0
	 ("00000000000000000000000000000000"),	 -- 1918	0
	 ("00000000000000000000000000000000"),	 -- 1917	0
	 ("00000000000000000000000000000000"),	 -- 1916	0
	 ("00000000000000000000000000000000"),	 -- 1915	0
	 ("00000000000000000000000000000000"),	 -- 1914	0
	 ("00000000000000000000000000000000"),	 -- 1913	0
	 ("00000000000000000000000000000000"),	 -- 1912	0
	 ("00000000000000000000000000000000"),	 -- 1911	0
	 ("00000000000000000000000000000000"),	 -- 1910	0
	 ("00000000000000000000000000000000"),	 -- 1909	0
	 ("00000000000000000000000000000000"),	 -- 1908	0
	 ("00000000000000000000000000000000"),	 -- 1907	0
	 ("00000000000000000000000000000000"),	 -- 1906	0
	 ("00000000000000000000000000000000"),	 -- 1905	0
	 ("00000000000000000000000000000000"),	 -- 1904	0
	 ("00000000000000000000000000000000"),	 -- 1903	0
	 ("00000000000000000000000000000000"),	 -- 1902	0
	 ("00000000000000000000000000000000"),	 -- 1901	0
	 ("00000000000000000000000000000000"),	 -- 1900	0
	 ("00000000000000000000000000000000"),	 -- 1899	0
	 ("00000000000000000000000000000000"),	 -- 1898	0
	 ("00000000000000000000000000000000"),	 -- 1897	0
	 ("00000000000000000000000000000000"),	 -- 1896	0
	 ("00000000000000000000000000000000"),	 -- 1895	0
	 ("00000000000000000000000000000000"),	 -- 1894	0
	 ("00000000000000000000000000000000"),	 -- 1893	0
	 ("00000000000000000000000000000000"),	 -- 1892	0
	 ("00000000000000000000000000000000"),	 -- 1891	0
	 ("00000000000000000000000000000000"),	 -- 1890	0
	 ("00000000000000000000000000000000"),	 -- 1889	0
	 ("00000000000000000000000000000000"),	 -- 1888	0
	 ("00000000000000000000000000000000"),	 -- 1887	0
	 ("00000000000000000000000000000000"),	 -- 1886	0
	 ("00000000000000000000000000000000"),	 -- 1885	0
	 ("00000000000000000000000000000000"),	 -- 1884	0
	 ("00000000000000000000000000000000"),	 -- 1883	0
	 ("00000000000000000000000000000000"),	 -- 1882	0
	 ("00000000000000000000000000000000"),	 -- 1881	0
	 ("00000000000000000000000000000000"),	 -- 1880	0
	 ("00000000000000000000000000000000"),	 -- 1879	0
	 ("00000000000000000000000000000000"),	 -- 1878	0
	 ("00000000000000000000000000000000"),	 -- 1877	0
	 ("00000000000000000000000000000000"),	 -- 1876	0
	 ("00000000000000000000000000000000"),	 -- 1875	0
	 ("00000000000000000000000000000000"),	 -- 1874	0
	 ("00000000000000000000000000000000"),	 -- 1873	0
	 ("00000000000000000000000000000000"),	 -- 1872	0
	 ("00000000000000000000000000000000"),	 -- 1871	0
	 ("00000000000000000000000000000000"),	 -- 1870	0
	 ("00000000000000000000000000000000"),	 -- 1869	0
	 ("00000000000000000000000000000000"),	 -- 1868	0
	 ("00000000000000000000000000000000"),	 -- 1867	0
	 ("00000000000000000000000000000000"),	 -- 1866	0
	 ("00000000000000000000000000000000"),	 -- 1865	0
	 ("00000000000000000000000000000000"),	 -- 1864	0
	 ("00000000000000000000000000000000"),	 -- 1863	0
	 ("00000000000000000000000000000000"),	 -- 1862	0
	 ("00000000000000000000000000000000"),	 -- 1861	0
	 ("00000000000000000000000000000000"),	 -- 1860	0
	 ("00000000000000000000000000000000"),	 -- 1859	0
	 ("00000000000000000000000000000000"),	 -- 1858	0
	 ("00000000000000000000000000000000"),	 -- 1857	0
	 ("00000000000000000000000000000000"),	 -- 1856	0
	 ("00000000000000000000000000000000"),	 -- 1855	0
	 ("00000000000000000000000000000000"),	 -- 1854	0
	 ("00000000000000000000000000000000"),	 -- 1853	0
	 ("00000000000000000000000000000000"),	 -- 1852	0
	 ("00000000000000000000000000000000"),	 -- 1851	0
	 ("00000000000000000000000000000000"),	 -- 1850	0
	 ("00000000000000000000000000000000"),	 -- 1849	0
	 ("00000000000000000000000000000000"),	 -- 1848	0
	 ("00000000000000000000000000000000"),	 -- 1847	0
	 ("00000000000000000000000000000000"),	 -- 1846	0
	 ("00000000000000000000000000000000"),	 -- 1845	0
	 ("00000000000000000000000000000000"),	 -- 1844	0
	 ("00000000000000000000000000000000"),	 -- 1843	0
	 ("00000000000000000000000000000000"),	 -- 1842	0
	 ("00000000000000000000000000000000"),	 -- 1841	0
	 ("00000000000000000000000000000000"),	 -- 1840	0
	 ("00000000000000000000000000000000"),	 -- 1839	0
	 ("00000000000000000000000000000000"),	 -- 1838	0
	 ("00000000000000000000000000000000"),	 -- 1837	0
	 ("00000000000000000000000000000000"),	 -- 1836	0
	 ("00000000000000000000000000000000"),	 -- 1835	0
	 ("00000000000000000000000000000000"),	 -- 1834	0
	 ("00000000000000000000000000000000"),	 -- 1833	0
	 ("00000000000000000000000000000000"),	 -- 1832	0
	 ("00000000000000000000000000000000"),	 -- 1831	0
	 ("00000000000000000000000000000000"),	 -- 1830	0
	 ("00000000000000000000000000000000"),	 -- 1829	0
	 ("00000000000000000000000000000000"),	 -- 1828	0
	 ("00000000000000000000000000000000"),	 -- 1827	0
	 ("00000000000000000000000000000000"),	 -- 1826	0
	 ("00000000000000000000000000000000"),	 -- 1825	0
	 ("00000000000000000000000000000000"),	 -- 1824	0
	 ("00000000000000000000000000000000"),	 -- 1823	0
	 ("00000000000000000000000000000000"),	 -- 1822	0
	 ("00000000000000000000000000000000"),	 -- 1821	0
	 ("00000000000000000000000000000000"),	 -- 1820	0
	 ("00000000000000000000000000000000"),	 -- 1819	0
	 ("00000000000000000000000000000000"),	 -- 1818	0
	 ("00000000000000000000000000000000"),	 -- 1817	0
	 ("00000000000000000000000000000000"),	 -- 1816	0
	 ("00000000000000000000000000000000"),	 -- 1815	0
	 ("00000000000000000000000000000000"),	 -- 1814	0
	 ("00000000000000000000000000000000"),	 -- 1813	0
	 ("00000000000000000000000000000000"),	 -- 1812	0
	 ("00000000000000000000000000000000"),	 -- 1811	0
	 ("00000000000000000000000000000000"),	 -- 1810	0
	 ("00000000000000000000000000000000"),	 -- 1809	0
	 ("00000000000000000000000000000000"),	 -- 1808	0
	 ("00000000000000000000000000000000"),	 -- 1807	0
	 ("00000000000000000000000000000000"),	 -- 1806	0
	 ("00000000000000000000000000000000"),	 -- 1805	0
	 ("00000000000000000000000000000000"),	 -- 1804	0
	 ("00000000000000000000000000000000"),	 -- 1803	0
	 ("00000000000000000000000000000000"),	 -- 1802	0
	 ("00000000000000000000000000000000"),	 -- 1801	0
	 ("00000000000000000000000000000000"),	 -- 1800	0
	 ("00000000000000000000000000000000"),	 -- 1799	0
	 ("00000000000000000000000000000000"),	 -- 1798	0
	 ("00000000000000000000000000000000"),	 -- 1797	0
	 ("00000000000000000000000000000000"),	 -- 1796	0
	 ("00000000000000000000000000000000"),	 -- 1795	0
	 ("00000000000000000000000000000000"),	 -- 1794	0
	 ("00000000000000000000000000000000"),	 -- 1793	0
	 ("00000000000000000000000000000000"),	 -- 1792	0
	 ("00000000000000000000000000000000"),	 -- 1791	0
	 ("00000000000000000000000000000000"),	 -- 1790	0
	 ("00000000000000000000000000000000"),	 -- 1789	0
	 ("00000000000000000000000000000000"),	 -- 1788	0
	 ("00000000000000000000000000000000"),	 -- 1787	0
	 ("00000000000000000000000000000000"),	 -- 1786	0
	 ("00000000000000000000000000000000"),	 -- 1785	0
	 ("00000000000000000000000000000000"),	 -- 1784	0
	 ("00000000000000000000000000000000"),	 -- 1783	0
	 ("00000000000000000000000000000000"),	 -- 1782	0
	 ("00000000000000000000000000000000"),	 -- 1781	0
	 ("00000000000000000000000000000000"),	 -- 1780	0
	 ("00000000000000000000000000000000"),	 -- 1779	0
	 ("00000000000000000000000000000000"),	 -- 1778	0
	 ("00000000000000000000000000000000"),	 -- 1777	0
	 ("00000000000000000000000000000000"),	 -- 1776	0
	 ("00000000000000000000000000000000"),	 -- 1775	0
	 ("00000000000000000000000000000000"),	 -- 1774	0
	 ("00000000000000000000000000000000"),	 -- 1773	0
	 ("00000000000000000000000000000000"),	 -- 1772	0
	 ("00000000000000000000000000000000"),	 -- 1771	0
	 ("00000000000000000000000000000000"),	 -- 1770	0
	 ("00000000000000000000000000000000"),	 -- 1769	0
	 ("00000000000000000000000000000000"),	 -- 1768	0
	 ("00000000000000000000000000000000"),	 -- 1767	0
	 ("00000000000000000000000000000000"),	 -- 1766	0
	 ("00000000000000000000000000000000"),	 -- 1765	0
	 ("00000000000000000000000000000000"),	 -- 1764	0
	 ("00000000000000000000000000000000"),	 -- 1763	0
	 ("00000000000000000000000000000000"),	 -- 1762	0
	 ("00000000000000000000000000000000"),	 -- 1761	0
	 ("00000000000000000000000000000000"),	 -- 1760	0
	 ("00000000000000000000000000000000"),	 -- 1759	0
	 ("00000000000000000000000000000000"),	 -- 1758	0
	 ("00000000000000000000000000000000"),	 -- 1757	0
	 ("00000000000000000000000000000000"),	 -- 1756	0
	 ("00000000000000000000000000000000"),	 -- 1755	0
	 ("00000000000000000000000000000000"),	 -- 1754	0
	 ("00000000000000000000000000000000"),	 -- 1753	0
	 ("00000000000000000000000000000000"),	 -- 1752	0
	 ("00000000000000000000000000000000"),	 -- 1751	0
	 ("00000000000000000000000000000000"),	 -- 1750	0
	 ("00000000000000000000000000000000"),	 -- 1749	0
	 ("00000000000000000000000000000000"),	 -- 1748	0
	 ("00000000000000000000000000000000"),	 -- 1747	0
	 ("00000000000000000000000000000000"),	 -- 1746	0
	 ("00000000000000000000000000000000"),	 -- 1745	0
	 ("00000000000000000000000000000000"),	 -- 1744	0
	 ("00000000000000000000000000000000"),	 -- 1743	0
	 ("00000000000000000000000000000000"),	 -- 1742	0
	 ("00000000000000000000000000000000"),	 -- 1741	0
	 ("00000000000000000000000000000000"),	 -- 1740	0
	 ("00000000000000000000000000000000"),	 -- 1739	0
	 ("00000000000000000000000000000000"),	 -- 1738	0
	 ("00000000000000000000000000000000"),	 -- 1737	0
	 ("00000000000000000000000000000000"),	 -- 1736	0
	 ("00000000000000000000000000000000"),	 -- 1735	0
	 ("00000000000000000000000000000000"),	 -- 1734	0
	 ("00000000000000000000000000000000"),	 -- 1733	0
	 ("00000000000000000000000000000000"),	 -- 1732	0
	 ("00000000000000000000000000000000"),	 -- 1731	0
	 ("00000000000000000000000000000000"),	 -- 1730	0
	 ("00000000000000000000000000000000"),	 -- 1729	0
	 ("00000000000000000000000000000000"),	 -- 1728	0
	 ("00000000000000000000000000000000"),	 -- 1727	0
	 ("00000000000000000000000000000000"),	 -- 1726	0
	 ("00000000000000000000000000000000"),	 -- 1725	0
	 ("00000000000000000000000000000000"),	 -- 1724	0
	 ("00000000000000000000000000000000"),	 -- 1723	0
	 ("00000000000000000000000000000000"),	 -- 1722	0
	 ("00000000000000000000000000000000"),	 -- 1721	0
	 ("00000000000000000000000000000000"),	 -- 1720	0
	 ("00000000000000000000000000000000"),	 -- 1719	0
	 ("00000000000000000000000000000000"),	 -- 1718	0
	 ("00000000000000000000000000000000"),	 -- 1717	0
	 ("00000000000000000000000000000000"),	 -- 1716	0
	 ("00000000000000000000000000000000"),	 -- 1715	0
	 ("00000000000000000000000000000000"),	 -- 1714	0
	 ("00000000000000000000000000000000"),	 -- 1713	0
	 ("00000000000000000000000000000000"),	 -- 1712	0
	 ("00000000000000000000000000000000"),	 -- 1711	0
	 ("00000000000000000000000000000000"),	 -- 1710	0
	 ("00000000000000000000000000000000"),	 -- 1709	0
	 ("00000000000000000000000000000000"),	 -- 1708	0
	 ("00000000000000000000000000000000"),	 -- 1707	0
	 ("00000000000000000000000000000000"),	 -- 1706	0
	 ("00000000000000000000000000000000"),	 -- 1705	0
	 ("00000000000000000000000000000000"),	 -- 1704	0
	 ("00000000000000000000000000000000"),	 -- 1703	0
	 ("00000000000000000000000000000000"),	 -- 1702	0
	 ("00000000000000000000000000000000"),	 -- 1701	0
	 ("00000000000000000000000000000000"),	 -- 1700	0
	 ("00000000000000000000000000000000"),	 -- 1699	0
	 ("00000000000000000000000000000000"),	 -- 1698	0
	 ("00000000000000000000000000000000"),	 -- 1697	0
	 ("00000000000000000000000000000000"),	 -- 1696	0
	 ("00000000000000000000000000000000"),	 -- 1695	0
	 ("00000000000000000000000000000000"),	 -- 1694	0
	 ("00000000000000000000000000000000"),	 -- 1693	0
	 ("00000000000000000000000000000000"),	 -- 1692	0
	 ("00000000000000000000000000000000"),	 -- 1691	0
	 ("00000000000000000000000000000000"),	 -- 1690	0
	 ("00000000000000000000000000000000"),	 -- 1689	0
	 ("00000000000000000000000000000000"),	 -- 1688	0
	 ("00000000000000000000000000000000"),	 -- 1687	0
	 ("00000000000000000000000000000000"),	 -- 1686	0
	 ("00000000000000000000000000000000"),	 -- 1685	0
	 ("00000000000000000000000000000000"),	 -- 1684	0
	 ("00000000000000000000000000000000"),	 -- 1683	0
	 ("00000000000000000000000000000000"),	 -- 1682	0
	 ("00000000000000000000000000000000"),	 -- 1681	0
	 ("00000000000000000000000000000000"),	 -- 1680	0
	 ("00000000000000000000000000000000"),	 -- 1679	0
	 ("00000000000000000000000000000000"),	 -- 1678	0
	 ("00000000000000000000000000000000"),	 -- 1677	0
	 ("00000000000000000000000000000000"),	 -- 1676	0
	 ("00000000000000000000000000000000"),	 -- 1675	0
	 ("00000000000000000000000000000000"),	 -- 1674	0
	 ("00000000000000000000000000000000"),	 -- 1673	0
	 ("00000000000000000000000000000000"),	 -- 1672	0
	 ("00000000000000000000000000000000"),	 -- 1671	0
	 ("00000000000000000000000000000000"),	 -- 1670	0
	 ("00000000000000000000000000000000"),	 -- 1669	0
	 ("00000000000000000000000000000000"),	 -- 1668	0
	 ("00000000000000000000000000000000"),	 -- 1667	0
	 ("00000000000000000000000000000000"),	 -- 1666	0
	 ("00000000000000000000000000000000"),	 -- 1665	0
	 ("00000000000000000000000000000000"),	 -- 1664	0
	 ("00000000000000000000000000000000"),	 -- 1663	0
	 ("00000000000000000000000000000000"),	 -- 1662	0
	 ("00000000000000000000000000000000"),	 -- 1661	0
	 ("00000000000000000000000000000000"),	 -- 1660	0
	 ("00000000000000000000000000000000"),	 -- 1659	0
	 ("00000000000000000000000000000000"),	 -- 1658	0
	 ("00000000000000000000000000000000"),	 -- 1657	0
	 ("00000000000000000000000000000000"),	 -- 1656	0
	 ("00000000000000000000000000000000"),	 -- 1655	0
	 ("00000000000000000000000000000000"),	 -- 1654	0
	 ("00000000000000000000000000000000"),	 -- 1653	0
	 ("00000000000000000000000000000000"),	 -- 1652	0
	 ("00000000000000000000000000000000"),	 -- 1651	0
	 ("00000000000000000000000000000000"),	 -- 1650	0
	 ("00000000000000000000000000000000"),	 -- 1649	0
	 ("00000000000000000000000000000000"),	 -- 1648	0
	 ("00000000000000000000000000000000"),	 -- 1647	0
	 ("00000000000000000000000000000000"),	 -- 1646	0
	 ("00000000000000000000000000000000"),	 -- 1645	0
	 ("00000000000000000000000000000000"),	 -- 1644	0
	 ("00000000000000000000000000000000"),	 -- 1643	0
	 ("00000000000000000000000000000000"),	 -- 1642	0
	 ("00000000000000000000000000000000"),	 -- 1641	0
	 ("00000000000000000000000000000000"),	 -- 1640	0
	 ("00000000000000000000000000000000"),	 -- 1639	0
	 ("00000000000000000000000000000000"),	 -- 1638	0
	 ("00000000000000000000000000000000"),	 -- 1637	0
	 ("00000000000000000000000000000000"),	 -- 1636	0
	 ("00000000000000000000000000000000"),	 -- 1635	0
	 ("00000000000000000000000000000000"),	 -- 1634	0
	 ("00000000000000000000000000000000"),	 -- 1633	0
	 ("00000000000000000000000000000000"),	 -- 1632	0
	 ("00000000000000000000000000000000"),	 -- 1631	0
	 ("00000000000000000000000000000000"),	 -- 1630	0
	 ("00000000000000000000000000000000"),	 -- 1629	0
	 ("00000000000000000000000000000000"),	 -- 1628	0
	 ("00000000000000000000000000000000"),	 -- 1627	0
	 ("00000000000000000000000000000000"),	 -- 1626	0
	 ("00000000000000000000000000000000"),	 -- 1625	0
	 ("00000000000000000000000000000000"),	 -- 1624	0
	 ("00000000000000000000000000000000"),	 -- 1623	0
	 ("00000000000000000000000000000000"),	 -- 1622	0
	 ("00000000000000000000000000000000"),	 -- 1621	0
	 ("00000000000000000000000000000000"),	 -- 1620	0
	 ("00000000000000000000000000000000"),	 -- 1619	0
	 ("00000000000000000000000000000000"),	 -- 1618	0
	 ("00000000000000000000000000000000"),	 -- 1617	0
	 ("00000000000000000000000000000000"),	 -- 1616	0
	 ("00000000000000000000000000000000"),	 -- 1615	0
	 ("00000000000000000000000000000000"),	 -- 1614	0
	 ("00000000000000000000000000000000"),	 -- 1613	0
	 ("00000000000000000000000000000000"),	 -- 1612	0
	 ("00000000000000000000000000000000"),	 -- 1611	0
	 ("00000000000000000000000000000000"),	 -- 1610	0
	 ("00000000000000000000000000000000"),	 -- 1609	0
	 ("00000000000000000000000000000000"),	 -- 1608	0
	 ("00000000000000000000000000000000"),	 -- 1607	0
	 ("00000000000000000000000000000000"),	 -- 1606	0
	 ("00000000000000000000000000000000"),	 -- 1605	0
	 ("00000000000000000000000000000000"),	 -- 1604	0
	 ("00000000000000000000000000000000"),	 -- 1603	0
	 ("00000000000000000000000000000000"),	 -- 1602	0
	 ("00000000000000000000000000000000"),	 -- 1601	0
	 ("00000000000000000000000000000000"),	 -- 1600	0
	 ("00000000000000000000000000000000"),	 -- 1599	0
	 ("00000000000000000000000000000000"),	 -- 1598	0
	 ("00000000000000000000000000000000"),	 -- 1597	0
	 ("00000000000000000000000000000000"),	 -- 1596	0
	 ("00000000000000000000000000000000"),	 -- 1595	0
	 ("00000000000000000000000000000000"),	 -- 1594	0
	 ("00000000000000000000000000000000"),	 -- 1593	0
	 ("00000000000000000000000000000000"),	 -- 1592	0
	 ("00000000000000000000000000000000"),	 -- 1591	0
	 ("00000000000000000000000000000000"),	 -- 1590	0
	 ("00000000000000000000000000000000"),	 -- 1589	0
	 ("00000000000000000000000000000000"),	 -- 1588	0
	 ("00000000000000000000000000000000"),	 -- 1587	0
	 ("00000000000000000000000000000000"),	 -- 1586	0
	 ("00000000000000000000000000000000"),	 -- 1585	0
	 ("00000000000000000000000000000000"),	 -- 1584	0
	 ("00000000000000000000000000000000"),	 -- 1583	0
	 ("00000000000000000000000000000000"),	 -- 1582	0
	 ("00000000000000000000000000000000"),	 -- 1581	0
	 ("00000000000000000000000000000000"),	 -- 1580	0
	 ("00000000000000000000000000000000"),	 -- 1579	0
	 ("00000000000000000000000000000000"),	 -- 1578	0
	 ("00000000000000000000000000000000"),	 -- 1577	0
	 ("00000000000000000000000000000000"),	 -- 1576	0
	 ("00000000000000000000000000000000"),	 -- 1575	0
	 ("00000000000000000000000000000000"),	 -- 1574	0
	 ("00000000000000000000000000000000"),	 -- 1573	0
	 ("00000000000000000000000000000000"),	 -- 1572	0
	 ("00000000000000000000000000000000"),	 -- 1571	0
	 ("00000000000000000000000000000000"),	 -- 1570	0
	 ("00000000000000000000000000000000"),	 -- 1569	0
	 ("00000000000000000000000000000000"),	 -- 1568	0
	 ("00000000000000000000000000000000"),	 -- 1567	0
	 ("00000000000000000000000000000000"),	 -- 1566	0
	 ("00000000000000000000000000000000"),	 -- 1565	0
	 ("00000000000000000000000000000000"),	 -- 1564	0
	 ("00000000000000000000000000000000"),	 -- 1563	0
	 ("00000000000000000000000000000000"),	 -- 1562	0
	 ("00000000000000000000000000000000"),	 -- 1561	0
	 ("00000000000000000000000000000000"),	 -- 1560	0
	 ("00000000000000000000000000000000"),	 -- 1559	0
	 ("00000000000000000000000000000000"),	 -- 1558	0
	 ("00000000000000000000000000000000"),	 -- 1557	0
	 ("00000000000000000000000000000000"),	 -- 1556	0
	 ("00000000000000000000000000000000"),	 -- 1555	0
	 ("00000000000000000000000000000000"),	 -- 1554	0
	 ("00000000000000000000000000000000"),	 -- 1553	0
	 ("00000000000000000000000000000000"),	 -- 1552	0
	 ("00000000000000000000000000000000"),	 -- 1551	0
	 ("00000000000000000000000000000000"),	 -- 1550	0
	 ("00000000000000000000000000000000"),	 -- 1549	0
	 ("00000000000000000000000000000000"),	 -- 1548	0
	 ("00000000000000000000000000000000"),	 -- 1547	0
	 ("00000000000000000000000000000000"),	 -- 1546	0
	 ("00000000000000000000000000000000"),	 -- 1545	0
	 ("00000000000000000000000000000000"),	 -- 1544	0
	 ("00000000000000000000000000000000"),	 -- 1543	0
	 ("00000000000000000000000000000000"),	 -- 1542	0
	 ("00000000000000000000000000000000"),	 -- 1541	0
	 ("00000000000000000000000000000000"),	 -- 1540	0
	 ("00000000000000000000000000000000"),	 -- 1539	0
	 ("00000000000000000000000000000000"),	 -- 1538	0
	 ("00000000000000000000000000000000"),	 -- 1537	0
	 ("00000000000000000000000000000000"),	 -- 1536	0
	 ("00000000000000000000000000000000"),	 -- 1535	0
	 ("00000000000000000000000000000000"),	 -- 1534	0
	 ("00000000000000000000000000000000"),	 -- 1533	0
	 ("00000000000000000000000000000000"),	 -- 1532	0
	 ("00000000000000000000000000000000"),	 -- 1531	0
	 ("00000000000000000000000000000000"),	 -- 1530	0
	 ("00000000000000000000000000000000"),	 -- 1529	0
	 ("00000000000000000000000000000000"),	 -- 1528	0
	 ("00000000000000000000000000000000"),	 -- 1527	0
	 ("00000000000000000000000000000000"),	 -- 1526	0
	 ("00000000000000000000000000000000"),	 -- 1525	0
	 ("00000000000000000000000000000000"),	 -- 1524	0
	 ("00000000000000000000000000000000"),	 -- 1523	0
	 ("00000000000000000000000000000000"),	 -- 1522	0
	 ("00000000000000000000000000000000"),	 -- 1521	0
	 ("00000000000000000000000000000000"),	 -- 1520	0
	 ("00000000000000000000000000000000"),	 -- 1519	0
	 ("00000000000000000000000000000000"),	 -- 1518	0
	 ("00000000000000000000000000000000"),	 -- 1517	0
	 ("00000000000000000000000000000000"),	 -- 1516	0
	 ("00000000000000000000000000000000"),	 -- 1515	0
	 ("00000000000000000000000000000000"),	 -- 1514	0
	 ("00000000000000000000000000000000"),	 -- 1513	0
	 ("00000000000000000000000000000000"),	 -- 1512	0
	 ("00000000000000000000000000000000"),	 -- 1511	0
	 ("00000000000000000000000000000000"),	 -- 1510	0
	 ("00000000000000000000000000000000"),	 -- 1509	0
	 ("00000000000000000000000000000000"),	 -- 1508	0
	 ("00000000000000000000000000000000"),	 -- 1507	0
	 ("00000000000000000000000000000000"),	 -- 1506	0
	 ("00000000000000000000000000000000"),	 -- 1505	0
	 ("00000000000000000000000000000000"),	 -- 1504	0
	 ("00000000000000000000000000000000"),	 -- 1503	0
	 ("00000000000000000000000000000000"),	 -- 1502	0
	 ("00000000000000000000000000000000"),	 -- 1501	0
	 ("00000000000000000000000000000000"),	 -- 1500	0
	 ("00000000000000000000000000000000"),	 -- 1499	0
	 ("00000000000000000000000000000000"),	 -- 1498	0
	 ("00000000000000000000000000000000"),	 -- 1497	0
	 ("00000000000000000000000000000000"),	 -- 1496	0
	 ("00000000000000000000000000000000"),	 -- 1495	0
	 ("00000000000000000000000000000000"),	 -- 1494	0
	 ("00000000000000000000000000000000"),	 -- 1493	0
	 ("00000000000000000000000000000000"),	 -- 1492	0
	 ("00000000000000000000000000000000"),	 -- 1491	0
	 ("00000000000000000000000000000000"),	 -- 1490	0
	 ("00000000000000000000000000000000"),	 -- 1489	0
	 ("00000000000000000000000000000000"),	 -- 1488	0
	 ("00000000000000000000000000000000"),	 -- 1487	0
	 ("00000000000000000000000000000000"),	 -- 1486	0
	 ("00000000000000000000000000000000"),	 -- 1485	0
	 ("00000000000000000000000000000000"),	 -- 1484	0
	 ("00000000000000000000000000000000"),	 -- 1483	0
	 ("00000000000000000000000000000000"),	 -- 1482	0
	 ("00000000000000000000000000000000"),	 -- 1481	0
	 ("00000000000000000000000000000000"),	 -- 1480	0
	 ("00000000000000000000000000000000"),	 -- 1479	0
	 ("00000000000000000000000000000000"),	 -- 1478	0
	 ("00000000000000000000000000000000"),	 -- 1477	0
	 ("00000000000000000000000000000000"),	 -- 1476	0
	 ("00000000000000000000000000000000"),	 -- 1475	0
	 ("00000000000000000000000000000000"),	 -- 1474	0
	 ("00000000000000000000000000000000"),	 -- 1473	0
	 ("00000000000000000000000000000000"),	 -- 1472	0
	 ("00000000000000000000000000000000"),	 -- 1471	0
	 ("00000000000000000000000000000000"),	 -- 1470	0
	 ("00000000000000000000000000000000"),	 -- 1469	0
	 ("00000000000000000000000000000000"),	 -- 1468	0
	 ("00000000000000000000000000000000"),	 -- 1467	0
	 ("00000000000000000000000000000000"),	 -- 1466	0
	 ("00000000000000000000000000000000"),	 -- 1465	0
	 ("00000000000000000000000000000000"),	 -- 1464	0
	 ("00000000000000000000000000000000"),	 -- 1463	0
	 ("00000000000000000000000000000000"),	 -- 1462	0
	 ("00000000000000000000000000000000"),	 -- 1461	0
	 ("00000000000000000000000000000000"),	 -- 1460	0
	 ("00000000000000000000000000000000"),	 -- 1459	0
	 ("00000000000000000000000000000000"),	 -- 1458	0
	 ("00000000000000000000000000000000"),	 -- 1457	0
	 ("00000000000000000000000000000000"),	 -- 1456	0
	 ("00000000000000000000000000000000"),	 -- 1455	0
	 ("00000000000000000000000000000000"),	 -- 1454	0
	 ("00000000000000000000000000000000"),	 -- 1453	0
	 ("00000000000000000000000000000000"),	 -- 1452	0
	 ("00000000000000000000000000000000"),	 -- 1451	0
	 ("00000000000000000000000000000000"),	 -- 1450	0
	 ("00000000000000000000000000000000"),	 -- 1449	0
	 ("00000000000000000000000000000000"),	 -- 1448	0
	 ("00000000000000000000000000000000"),	 -- 1447	0
	 ("00000000000000000000000000000000"),	 -- 1446	0
	 ("00000000000000000000000000000000"),	 -- 1445	0
	 ("00000000000000000000000000000000"),	 -- 1444	0
	 ("00000000000000000000000000000000"),	 -- 1443	0
	 ("00000000000000000000000000000000"),	 -- 1442	0
	 ("00000000000000000000000000000000"),	 -- 1441	0
	 ("00000000000000000000000000000000"),	 -- 1440	0
	 ("00000000000000000000000000000000"),	 -- 1439	0
	 ("00000000000000000000000000000000"),	 -- 1438	0
	 ("00000000000000000000000000000000"),	 -- 1437	0
	 ("00000000000000000000000000000000"),	 -- 1436	0
	 ("00000000000000000000000000000000"),	 -- 1435	0
	 ("00000000000000000000000000000000"),	 -- 1434	0
	 ("00000000000000000000000000000000"),	 -- 1433	0
	 ("00000000000000000000000000000000"),	 -- 1432	0
	 ("00000000000000000000000000000000"),	 -- 1431	0
	 ("00000000000000000000000000000000"),	 -- 1430	0
	 ("00000000000000000000000000000000"),	 -- 1429	0
	 ("00000000000000000000000000000000"),	 -- 1428	0
	 ("00000000000000000000000000000000"),	 -- 1427	0
	 ("00000000000000000000000000000000"),	 -- 1426	0
	 ("00000000000000000000000000000000"),	 -- 1425	0
	 ("00000000000000000000000000000000"),	 -- 1424	0
	 ("00000000000000000000000000000000"),	 -- 1423	0
	 ("00000000000000000000000000000000"),	 -- 1422	0
	 ("00000000000000000000000000000000"),	 -- 1421	0
	 ("00000000000000000000000000000000"),	 -- 1420	0
	 ("00000000000000000000000000000000"),	 -- 1419	0
	 ("00000000000000000000000000000000"),	 -- 1418	0
	 ("00000000000000000000000000000000"),	 -- 1417	0
	 ("00000000000000000000000000000000"),	 -- 1416	0
	 ("00000000000000000000000000000000"),	 -- 1415	0
	 ("00000000000000000000000000000000"),	 -- 1414	0
	 ("00000000000000000000000000000000"),	 -- 1413	0
	 ("00000000000000000000000000000000"),	 -- 1412	0
	 ("00000000000000000000000000000000"),	 -- 1411	0
	 ("00000000000000000000000000000000"),	 -- 1410	0
	 ("00000000000000000000000000000000"),	 -- 1409	0
	 ("00000000000000000000000000000000"),	 -- 1408	0
	 ("00000000000000000000000000000000"),	 -- 1407	0
	 ("00000000000000000000000000000000"),	 -- 1406	0
	 ("00000000000000000000000000000000"),	 -- 1405	0
	 ("00000000000000000000000000000000"),	 -- 1404	0
	 ("00000000000000000000000000000000"),	 -- 1403	0
	 ("00000000000000000000000000000000"),	 -- 1402	0
	 ("00000000000000000000000000000000"),	 -- 1401	0
	 ("00000000000000000000000000000000"),	 -- 1400	0
	 ("00000000000000000000000000000000"),	 -- 1399	0
	 ("00000000000000000000000000000000"),	 -- 1398	0
	 ("00000000000000000000000000000000"),	 -- 1397	0
	 ("00000000000000000000000000000000"),	 -- 1396	0
	 ("00000000000000000000000000000000"),	 -- 1395	0
	 ("00000000000000000000000000000000"),	 -- 1394	0
	 ("00000000000000000000000000000000"),	 -- 1393	0
	 ("00000000000000000000000000000000"),	 -- 1392	0
	 ("00000000000000000000000000000000"),	 -- 1391	0
	 ("00000000000000000000000000000000"),	 -- 1390	0
	 ("00000000000000000000000000000000"),	 -- 1389	0
	 ("00000000000000000000000000000000"),	 -- 1388	0
	 ("00000000000000000000000000000000"),	 -- 1387	0
	 ("00000000000000000000000000000000"),	 -- 1386	0
	 ("00000000000000000000000000000000"),	 -- 1385	0
	 ("00000000000000000000000000000000"),	 -- 1384	0
	 ("00000000000000000000000000000000"),	 -- 1383	0
	 ("00000000000000000000000000000000"),	 -- 1382	0
	 ("00000000000000000000000000000000"),	 -- 1381	0
	 ("00000000000000000000000000000000"),	 -- 1380	0
	 ("00000000000000000000000000000000"),	 -- 1379	0
	 ("00000000000000000000000000000000"),	 -- 1378	0
	 ("00000000000000000000000000000000"),	 -- 1377	0
	 ("00000000000000000000000000000000"),	 -- 1376	0
	 ("00000000000000000000000000000000"),	 -- 1375	0
	 ("00000000000000000000000000000000"),	 -- 1374	0
	 ("00000000000000000000000000000000"),	 -- 1373	0
	 ("00000000000000000000000000000000"),	 -- 1372	0
	 ("00000000000000000000000000000000"),	 -- 1371	0
	 ("00000000000000000000000000000000"),	 -- 1370	0
	 ("00000000000000000000000000000000"),	 -- 1369	0
	 ("00000000000000000000000000000000"),	 -- 1368	0
	 ("00000000000000000000000000000000"),	 -- 1367	0
	 ("00000000000000000000000000000000"),	 -- 1366	0
	 ("00000000000000000000000000000000"),	 -- 1365	0
	 ("00000000000000000000000000000000"),	 -- 1364	0
	 ("00000000000000000000000000000000"),	 -- 1363	0
	 ("00000000000000000000000000000000"),	 -- 1362	0
	 ("00000000000000000000000000000000"),	 -- 1361	0
	 ("00000000000000000000000000000000"),	 -- 1360	0
	 ("00000000000000000000000000000000"),	 -- 1359	0
	 ("00000000000000000000000000000000"),	 -- 1358	0
	 ("00000000000000000000000000000000"),	 -- 1357	0
	 ("00000000000000000000000000000000"),	 -- 1356	0
	 ("00000000000000000000000000000000"),	 -- 1355	0
	 ("00000000000000000000000000000000"),	 -- 1354	0
	 ("00000000000000000000000000000000"),	 -- 1353	0
	 ("00000000000000000000000000000000"),	 -- 1352	0
	 ("00000000000000000000000000000000"),	 -- 1351	0
	 ("00000000000000000000000000000000"),	 -- 1350	0
	 ("00000000000000000000000000000000"),	 -- 1349	0
	 ("00000000000000000000000000000000"),	 -- 1348	0
	 ("00000000000000000000000000000000"),	 -- 1347	0
	 ("00000000000000000000000000000000"),	 -- 1346	0
	 ("00000000000000000000000000000000"),	 -- 1345	0
	 ("00000000000000000000000000000000"),	 -- 1344	0
	 ("00000000000000000000000000000000"),	 -- 1343	0
	 ("00000000000000000000000000000000"),	 -- 1342	0
	 ("00000000000000000000000000000000"),	 -- 1341	0
	 ("00000000000000000000000000000000"),	 -- 1340	0
	 ("00000000000000000000000000000000"),	 -- 1339	0
	 ("00000000000000000000000000000000"),	 -- 1338	0
	 ("00000000000000000000000000000000"),	 -- 1337	0
	 ("00000000000000000000000000000000"),	 -- 1336	0
	 ("00000000000000000000000000000000"),	 -- 1335	0
	 ("00000000000000000000000000000000"),	 -- 1334	0
	 ("00000000000000000000000000000000"),	 -- 1333	0
	 ("00000000000000000000000000000000"),	 -- 1332	0
	 ("00000000000000000000000000000000"),	 -- 1331	0
	 ("00000000000000000000000000000000"),	 -- 1330	0
	 ("00000000000000000000000000000000"),	 -- 1329	0
	 ("00000000000000000000000000000000"),	 -- 1328	0
	 ("00000000000000000000000000000000"),	 -- 1327	0
	 ("00000000000000000000000000000000"),	 -- 1326	0
	 ("00000000000000000000000000000000"),	 -- 1325	0
	 ("00000000000000000000000000000000"),	 -- 1324	0
	 ("00000000000000000000000000000000"),	 -- 1323	0
	 ("00000000000000000000000000000000"),	 -- 1322	0
	 ("00000000000000000000000000000000"),	 -- 1321	0
	 ("00000000000000000000000000000000"),	 -- 1320	0
	 ("00000000000000000000000000000000"),	 -- 1319	0
	 ("00000000000000000000000000000000"),	 -- 1318	0
	 ("00000000000000000000000000000000"),	 -- 1317	0
	 ("00000000000000000000000000000000"),	 -- 1316	0
	 ("00000000000000000000000000000000"),	 -- 1315	0
	 ("00000000000000000000000000000000"),	 -- 1314	0
	 ("00000000000000000000000000000000"),	 -- 1313	0
	 ("00000000000000000000000000000000"),	 -- 1312	0
	 ("00000000000000000000000000000000"),	 -- 1311	0
	 ("00000000000000000000000000000000"),	 -- 1310	0
	 ("00000000000000000000000000000000"),	 -- 1309	0
	 ("00000000000000000000000000000000"),	 -- 1308	0
	 ("00000000000000000000000000000000"),	 -- 1307	0
	 ("00000000000000000000000000000000"),	 -- 1306	0
	 ("00000000000000000000000000000000"),	 -- 1305	0
	 ("00000000000000000000000000000000"),	 -- 1304	0
	 ("00000000000000000000000000000000"),	 -- 1303	0
	 ("00000000000000000000000000000000"),	 -- 1302	0
	 ("00000000000000000000000000000000"),	 -- 1301	0
	 ("00000000000000000000000000000000"),	 -- 1300	0
	 ("00000000000000000000000000000000"),	 -- 1299	0
	 ("00000000000000000000000000000000"),	 -- 1298	0
	 ("00000000000000000000000000000000"),	 -- 1297	0
	 ("00000000000000000000000000000000"),	 -- 1296	0
	 ("00000000000000000000000000000000"),	 -- 1295	0
	 ("00000000000000000000000000000000"),	 -- 1294	0
	 ("00000000000000000000000000000000"),	 -- 1293	0
	 ("00000000000000000000000000000000"),	 -- 1292	0
	 ("00000000000000000000000000000000"),	 -- 1291	0
	 ("00000000000000000000000000000000"),	 -- 1290	0
	 ("00000000000000000000000000000000"),	 -- 1289	0
	 ("00000000000000000000000000000000"),	 -- 1288	0
	 ("00000000000000000000000000000000"),	 -- 1287	0
	 ("00000000000000000000000000000000"),	 -- 1286	0
	 ("00000000000000000000000000000000"),	 -- 1285	0
	 ("00000000000000000000000000000000"),	 -- 1284	0
	 ("00000000000000000000000000000000"),	 -- 1283	0
	 ("00000000000000000000000000000000"),	 -- 1282	0
	 ("00000000000000000000000000000000"),	 -- 1281	0
	 ("00000000000000000000000000000000"),	 -- 1280	0
	 ("00000000000000000000000000000000"),	 -- 1279	0
	 ("00000000000000000000000000000000"),	 -- 1278	0
	 ("00000000000000000000000000000000"),	 -- 1277	0
	 ("00000000000000000000000000000000"),	 -- 1276	0
	 ("00000000000000000000000000000000"),	 -- 1275	0
	 ("00000000000000000000000000000000"),	 -- 1274	0
	 ("00000000000000000000000000000000"),	 -- 1273	0
	 ("00000000000000000000000000000000"),	 -- 1272	0
	 ("00000000000000000000000000000000"),	 -- 1271	0
	 ("00000000000000000000000000000000"),	 -- 1270	0
	 ("00000000000000000000000000000000"),	 -- 1269	0
	 ("00000000000000000000000000000000"),	 -- 1268	0
	 ("00000000000000000000000000000000"),	 -- 1267	0
	 ("00000000000000000000000000000000"),	 -- 1266	0
	 ("00000000000000000000000000000000"),	 -- 1265	0
	 ("00000000000000000000000000000000"),	 -- 1264	0
	 ("00000000000000000000000000000000"),	 -- 1263	0
	 ("00000000000000000000000000000000"),	 -- 1262	0
	 ("00000000000000000000000000000000"),	 -- 1261	0
	 ("00000000000000000000000000000000"),	 -- 1260	0
	 ("00000000000000000000000000000000"),	 -- 1259	0
	 ("00000000000000000000000000000000"),	 -- 1258	0
	 ("00000000000000000000000000000000"),	 -- 1257	0
	 ("00000000000000000000000000000000"),	 -- 1256	0
	 ("00000000000000000000000000000000"),	 -- 1255	0
	 ("00000000000000000000000000000000"),	 -- 1254	0
	 ("00000000000000000000000000000000"),	 -- 1253	0
	 ("00000000000000000000000000000000"),	 -- 1252	0
	 ("00000000000000000000000000000000"),	 -- 1251	0
	 ("00000000000000000000000000000000"),	 -- 1250	0
	 ("00000000000000000000000000000000"),	 -- 1249	0
	 ("00000000000000000000000000000000"),	 -- 1248	0
	 ("00000000000000000000000000000000"),	 -- 1247	0
	 ("00000000000000000000000000000000"),	 -- 1246	0
	 ("00000000000000000000000000000000"),	 -- 1245	0
	 ("00000000000000000000000000000000"),	 -- 1244	0
	 ("00000000000000000000000000000000"),	 -- 1243	0
	 ("00000000000000000000000000000000"),	 -- 1242	0
	 ("00000000000000000000000000000000"),	 -- 1241	0
	 ("00000000000000000000000000000000"),	 -- 1240	0
	 ("00000000000000000000000000000000"),	 -- 1239	0
	 ("00000000000000000000000000000000"),	 -- 1238	0
	 ("00000000000000000000000000000000"),	 -- 1237	0
	 ("00000000000000000000000000000000"),	 -- 1236	0
	 ("00000000000000000000000000000000"),	 -- 1235	0
	 ("00000000000000000000000000000000"),	 -- 1234	0
	 ("00000000000000000000000000000000"),	 -- 1233	0
	 ("00000000000000000000000000000000"),	 -- 1232	0
	 ("00000000000000000000000000000000"),	 -- 1231	0
	 ("00000000000000000000000000000000"),	 -- 1230	0
	 ("00000000000000000000000000000000"),	 -- 1229	0
	 ("00000000000000000000000000000000"),	 -- 1228	0
	 ("00000000000000000000000000000000"),	 -- 1227	0
	 ("00000000000000000000000000000000"),	 -- 1226	0
	 ("00000000000000000000000000000000"),	 -- 1225	0
	 ("00000000000000000000000000000000"),	 -- 1224	0
	 ("00000000000000000000000000000000"),	 -- 1223	0
	 ("00000000000000000000000000000000"),	 -- 1222	0
	 ("00000000000000000000000000000000"),	 -- 1221	0
	 ("00000000000000000000000000000000"),	 -- 1220	0
	 ("00000000000000000000000000000000"),	 -- 1219	0
	 ("00000000000000000000000000000000"),	 -- 1218	0
	 ("00000000000000000000000000000000"),	 -- 1217	0
	 ("00000000000000000000000000000000"),	 -- 1216	0
	 ("00000000000000000000000000000000"),	 -- 1215	0
	 ("00000000000000000000000000000000"),	 -- 1214	0
	 ("00000000000000000000000000000000"),	 -- 1213	0
	 ("00000000000000000000000000000000"),	 -- 1212	0
	 ("00000000000000000000000000000000"),	 -- 1211	0
	 ("00000000000000000000000000000000"),	 -- 1210	0
	 ("00000000000000000000000000000000"),	 -- 1209	0
	 ("00000000000000000000000000000000"),	 -- 1208	0
	 ("00000000000000000000000000000000"),	 -- 1207	0
	 ("00000000000000000000000000000000"),	 -- 1206	0
	 ("00000000000000000000000000000000"),	 -- 1205	0
	 ("00000000000000000000000000000000"),	 -- 1204	0
	 ("00000000000000000000000000000000"),	 -- 1203	0
	 ("00000000000000000000000000000000"),	 -- 1202	0
	 ("00000000000000000000000000000000"),	 -- 1201	0
	 ("00000000000000000000000000000000"),	 -- 1200	0
	 ("00000000000000000000000000000000"),	 -- 1199	0
	 ("00000000000000000000000000000000"),	 -- 1198	0
	 ("00000000000000000000000000000000"),	 -- 1197	0
	 ("00000000000000000000000000000000"),	 -- 1196	0
	 ("00000000000000000000000000000000"),	 -- 1195	0
	 ("00000000000000000000000000000000"),	 -- 1194	0
	 ("00000000000000000000000000000000"),	 -- 1193	0
	 ("00000000000000000000000000000000"),	 -- 1192	0
	 ("00000000000000000000000000000000"),	 -- 1191	0
	 ("00000000000000000000000000000000"),	 -- 1190	0
	 ("00000000000000000000000000000000"),	 -- 1189	0
	 ("00000000000000000000000000000000"),	 -- 1188	0
	 ("00000000000000000000000000000000"),	 -- 1187	0
	 ("00000000000000000000000000000000"),	 -- 1186	0
	 ("00000000000000000000000000000000"),	 -- 1185	0
	 ("00000000000000000000000000000000"),	 -- 1184	0
	 ("00000000000000000000000000000000"),	 -- 1183	0
	 ("00000000000000000000000000000000"),	 -- 1182	0
	 ("00000000000000000000000000000000"),	 -- 1181	0
	 ("00000000000000000000000000000000"),	 -- 1180	0
	 ("00000000000000000000000000000000"),	 -- 1179	0
	 ("00000000000000000000000000000000"),	 -- 1178	0
	 ("00000000000000000000000000000000"),	 -- 1177	0
	 ("00000000000000000000000000000000"),	 -- 1176	0
	 ("00000000000000000000000000000000"),	 -- 1175	0
	 ("00000000000000000000000000000000"),	 -- 1174	0
	 ("00000000000000000000000000000000"),	 -- 1173	0
	 ("00000000000000000000000000000000"),	 -- 1172	0
	 ("00000000000000000000000000000000"),	 -- 1171	0
	 ("00000000000000000000000000000000"),	 -- 1170	0
	 ("00000000000000000000000000000000"),	 -- 1169	0
	 ("00000000000000000000000000000000"),	 -- 1168	0
	 ("00000000000000000000000000000000"),	 -- 1167	0
	 ("00000000000000000000000000000000"),	 -- 1166	0
	 ("00000000000000000000000000000000"),	 -- 1165	0
	 ("00000000000000000000000000000000"),	 -- 1164	0
	 ("00000000000000000000000000000000"),	 -- 1163	0
	 ("00000000000000000000000000000000"),	 -- 1162	0
	 ("00000000000000000000000000000000"),	 -- 1161	0
	 ("00000000000000000000000000000000"),	 -- 1160	0
	 ("00000000000000000000000000000000"),	 -- 1159	0
	 ("00000000000000000000000000000000"),	 -- 1158	0
	 ("00000000000000000000000000000000"),	 -- 1157	0
	 ("00000000000000000000000000000000"),	 -- 1156	0
	 ("00000000000000000000000000000000"),	 -- 1155	0
	 ("00000000000000000000000000000000"),	 -- 1154	0
	 ("00000000000000000000000000000000"),	 -- 1153	0
	 ("00000000000000000000000000000000"),	 -- 1152	0
	 ("00000000000000000000000000000000"),	 -- 1151	0
	 ("00000000000000000000000000000000"),	 -- 1150	0
	 ("00000000000000000000000000000000"),	 -- 1149	0
	 ("00000000000000000000000000000000"),	 -- 1148	0
	 ("00000000000000000000000000000000"),	 -- 1147	0
	 ("00000000000000000000000000000000"),	 -- 1146	0
	 ("00000000000000000000000000000000"),	 -- 1145	0
	 ("00000000000000000000000000000000"),	 -- 1144	0
	 ("00000000000000000000000000000000"),	 -- 1143	0
	 ("00000000000000000000000000000000"),	 -- 1142	0
	 ("00000000000000000000000000000000"),	 -- 1141	0
	 ("00000000000000000000000000000000"),	 -- 1140	0
	 ("00000000000000000000000000000000"),	 -- 1139	0
	 ("00000000000000000000000000000000"),	 -- 1138	0
	 ("00000000000000000000000000000000"),	 -- 1137	0
	 ("00000000000000000000000000000000"),	 -- 1136	0
	 ("00000000000000000000000000000000"),	 -- 1135	0
	 ("00000000000000000000000000000000"),	 -- 1134	0
	 ("00000000000000000000000000000000"),	 -- 1133	0
	 ("00000000000000000000000000000000"),	 -- 1132	0
	 ("00000000000000000000000000000000"),	 -- 1131	0
	 ("00000000000000000000000000000000"),	 -- 1130	0
	 ("00000000000000000000000000000000"),	 -- 1129	0
	 ("00000000000000000000000000000000"),	 -- 1128	0
	 ("00000000000000000000000000000000"),	 -- 1127	0
	 ("00000000000000000000000000000000"),	 -- 1126	0
	 ("00000000000000000000000000000000"),	 -- 1125	0
	 ("00000000000000000000000000000000"),	 -- 1124	0
	 ("00000000000000000000000000000000"),	 -- 1123	0
	 ("00000000000000000000000000000000"),	 -- 1122	0
	 ("00000000000000000000000000000000"),	 -- 1121	0
	 ("00000000000000000000000000000000"),	 -- 1120	0
	 ("00000000000000000000000000000000"),	 -- 1119	0
	 ("00000000000000000000000000000000"),	 -- 1118	0
	 ("00000000000000000000000000000000"),	 -- 1117	0
	 ("00000000000000000000000000000000"),	 -- 1116	0
	 ("00000000000000000000000000000000"),	 -- 1115	0
	 ("00000000000000000000000000000000"),	 -- 1114	0
	 ("00000000000000000000000000000000"),	 -- 1113	0
	 ("00000000000000000000000000000000"),	 -- 1112	0
	 ("00000000000000000000000000000000"),	 -- 1111	0
	 ("00000000000000000000000000000000"),	 -- 1110	0
	 ("00000000000000000000000000000000"),	 -- 1109	0
	 ("00000000000000000000000000000000"),	 -- 1108	0
	 ("00000000000000000000000000000000"),	 -- 1107	0
	 ("00000000000000000000000000000000"),	 -- 1106	0
	 ("00000000000000000000000000000000"),	 -- 1105	0
	 ("00000000000000000000000000000000"),	 -- 1104	0
	 ("00000000000000000000000000000000"),	 -- 1103	0
	 ("00000000000000000000000000000000"),	 -- 1102	0
	 ("00000000000000000000000000000000"),	 -- 1101	0
	 ("00000000000000000000000000000000"),	 -- 1100	0
	 ("00000000000000000000000000000000"),	 -- 1099	0
	 ("00000000000000000000000000000000"),	 -- 1098	0
	 ("00000000000000000000000000000000"),	 -- 1097	0
	 ("00000000000000000000000000000000"),	 -- 1096	0
	 ("00000000000000000000000000000000"),	 -- 1095	0
	 ("00000000000000000000000000000000"),	 -- 1094	0
	 ("00000000000000000000000000000000"),	 -- 1093	0
	 ("00000000000000000000000000000000"),	 -- 1092	0
	 ("00000000000000000000000000000000"),	 -- 1091	0
	 ("00000000000000000000000000000000"),	 -- 1090	0
	 ("00000000000000000000000000000000"),	 -- 1089	0
	 ("00000000000000000000000000000000"),	 -- 1088	0
	 ("00000000000000000000000000000000"),	 -- 1087	0
	 ("00000000000000000000000000000000"),	 -- 1086	0
	 ("00000000000000000000000000000000"),	 -- 1085	0
	 ("00000000000000000000000000000000"),	 -- 1084	0
	 ("00000000000000000000000000000000"),	 -- 1083	0
	 ("00000000000000000000000000000000"),	 -- 1082	0
	 ("00000000000000000000000000000000"),	 -- 1081	0
	 ("00000000000000000000000000000000"),	 -- 1080	0
	 ("00000000000000000000000000000000"),	 -- 1079	0
	 ("00000000000000000000000000000000"),	 -- 1078	0
	 ("00000000000000000000000000000000"),	 -- 1077	0
	 ("00000000000000000000000000000000"),	 -- 1076	0
	 ("00000000000000000000000000000000"),	 -- 1075	0
	 ("00000000000000000000000000000000"),	 -- 1074	0
	 ("00000000000000000000000000000000"),	 -- 1073	0
	 ("00000000000000000000000000000000"),	 -- 1072	0
	 ("00000000000000000000000000000000"),	 -- 1071	0
	 ("00000000000000000000000000000000"),	 -- 1070	0
	 ("00000000000000000000000000000000"),	 -- 1069	0
	 ("00000000000000000000000000000000"),	 -- 1068	0
	 ("00000000000000000000000000000000"),	 -- 1067	0
	 ("00000000000000000000000000000000"),	 -- 1066	0
	 ("00000000000000000000000000000000"),	 -- 1065	0
	 ("00000000000000000000000000000000"),	 -- 1064	0
	 ("00000000000000000000000000000000"),	 -- 1063	0
	 ("00000000000000000000000000000000"),	 -- 1062	0
	 ("00000000000000000000000000000000"),	 -- 1061	0
	 ("00000000000000000000000000000000"),	 -- 1060	0
	 ("00000000000000000000000000000000"),	 -- 1059	0
	 ("00000000000000000000000000000000"),	 -- 1058	0
	 ("00000000000000000000000000000000"),	 -- 1057	0
	 ("00000000000000000000000000000000"),	 -- 1056	0
	 ("00000000000000000000000000000000"),	 -- 1055	0
	 ("00000000000000000000000000000000"),	 -- 1054	0
	 ("00000000000000000000000000000000"),	 -- 1053	0
	 ("00000000000000000000000000000000"),	 -- 1052	0
	 ("00000000000000000000000000000000"),	 -- 1051	0
	 ("00000000000000000000000000000000"),	 -- 1050	0
	 ("00000000000000000000000000000000"),	 -- 1049	0
	 ("00000000000000000000000000000000"),	 -- 1048	0
	 ("00000000000000000000000000000000"),	 -- 1047	0
	 ("00000000000000000000000000000000"),	 -- 1046	0
	 ("00000000000000000000000000000000"),	 -- 1045	0
	 ("00000000000000000000000000000000"),	 -- 1044	0
	 ("00000000000000000000000000000000"),	 -- 1043	0
	 ("00000000000000000000000000000000"),	 -- 1042	0
	 ("00000000000000000000000000000000"),	 -- 1041	0
	 ("00000000000000000000000000000000"),	 -- 1040	0
	 ("00000000000000000000000000000000"),	 -- 1039	0
	 ("00000000000000000000000000000000"),	 -- 1038	0
	 ("00000000000000000000000000000000"),	 -- 1037	0
	 ("00000000000000000000000000000000"),	 -- 1036	0
	 ("00000000000000000000000000000000"),	 -- 1035	0
	 ("00000000000000000000000000000000"),	 -- 1034	0
	 ("00000000000000000000000000000000"),	 -- 1033	0
	 ("00000000000000000000000000000000"),	 -- 1032	0
	 ("00000000000000000000000000000000"),	 -- 1031	0
	 ("00000000000000000000000000000000"),	 -- 1030	0
	 ("00000000000000000000000000000000"),	 -- 1029	0
	 ("00000000000000000000000000000000"),	 -- 1028	0
	 ("00000000000000000000000000000000"),	 -- 1027	0
	 ("00000000000000000000000000000000"),	 -- 1026	0
	 ("00000000000000000000000000000000"),	 -- 1025	0
	 ("00000000000000000000000000000000"),	 -- 1024	0
	 ("00000000000000000000000000000000"),	 -- 1023	0
	 ("00000000000000000000000000000000"),	 -- 1022	0
	 ("00000000000000000000000000000000"),	 -- 1021	0
	 ("00000000000000000000000000000000"),	 -- 1020	0
	 ("00000000000000000000000000000000"),	 -- 1019	0
	 ("00000000000000000000000000000000"),	 -- 1018	0
	 ("00000000000000000000000000000000"),	 -- 1017	0
	 ("00000000000000000000000000000000"),	 -- 1016	0
	 ("00000000000000000000000000000000"),	 -- 1015	0
	 ("00000000000000000000000000000000"),	 -- 1014	0
	 ("00000000000000000000000000000000"),	 -- 1013	0
	 ("00000000000000000000000000000000"),	 -- 1012	0
	 ("00000000000000000000000000000000"),	 -- 1011	0
	 ("00000000000000000000000000000000"),	 -- 1010	0
	 ("00000000000000000000000000000000"),	 -- 1009	0
	 ("00000000000000000000000000000000"),	 -- 1008	0
	 ("00000000000000000000000000000000"),	 -- 1007	0
	 ("00000000000000000000000000000000"),	 -- 1006	0
	 ("00000000000000000000000000000000"),	 -- 1005	0
	 ("00000000000000000000000000000000"),	 -- 1004	0
	 ("00000000000000000000000000000000"),	 -- 1003	0
	 ("00000000000000000000000000000000"),	 -- 1002	0
	 ("00000000000000000000000000000000"),	 -- 1001	0
	 ("00000000000000000000000000000000"),	 -- 1000	0
	 ("00000000000000000000000000000000"),	 -- 999	0
	 ("00000000000000000000000000000000"),	 -- 998	0
	 ("00000000000000000000000000000000"),	 -- 997	0
	 ("00000000000000000000000000000000"),	 -- 996	0
	 ("00000000000000000000000000000000"),	 -- 995	0
	 ("00000000000000000000000000000000"),	 -- 994	0
	 ("00000000000000000000000000000000"),	 -- 993	0
	 ("00000000000000000000000000000000"),	 -- 992	0
	 ("00000000000000000000000000000000"),	 -- 991	0
	 ("00000000000000000000000000000000"),	 -- 990	0
	 ("00000000000000000000000000000000"),	 -- 989	0
	 ("00000000000000000000000000000000"),	 -- 988	0
	 ("00000000000000000000000000000000"),	 -- 987	0
	 ("00000000000000000000000000000000"),	 -- 986	0
	 ("00000000000000000000000000000000"),	 -- 985	0
	 ("00000000000000000000000000000000"),	 -- 984	0
	 ("00000000000000000000000000000000"),	 -- 983	0
	 ("00000000000000000000000000000000"),	 -- 982	0
	 ("00000000000000000000000000000000"),	 -- 981	0
	 ("00000000000000000000000000000000"),	 -- 980	0
	 ("00000000000000000000000000000000"),	 -- 979	0
	 ("00000000000000000000000000000000"),	 -- 978	0
	 ("00000000000000000000000000000000"),	 -- 977	0
	 ("00000000000000000000000000000000"),	 -- 976	0
	 ("00000000000000000000000000000000"),	 -- 975	0
	 ("00000000000000000000000000000000"),	 -- 974	0
	 ("00000000000000000000000000000000"),	 -- 973	0
	 ("00000000000000000000000000000000"),	 -- 972	0
	 ("00000000000000000000000000000000"),	 -- 971	0
	 ("00000000000000000000000000000000"),	 -- 970	0
	 ("00000000000000000000000000000000"),	 -- 969	0
	 ("00000000000000000000000000000000"),	 -- 968	0
	 ("00000000000000000000000000000000"),	 -- 967	0
	 ("00000000000000000000000000000000"),	 -- 966	0
	 ("00000000000000000000000000000000"),	 -- 965	0
	 ("00000000000000000000000000000000"),	 -- 964	0
	 ("00000000000000000000000000000000"),	 -- 963	0
	 ("00000000000000000000000000000000"),	 -- 962	0
	 ("00000000000000000000000000000000"),	 -- 961	0
	 ("00000000000000000000000000000000"),	 -- 960	0
	 ("00000000000000000000000000000000"),	 -- 959	0
	 ("00000000000000000000000000000000"),	 -- 958	0
	 ("00000000000000000000000000000000"),	 -- 957	0
	 ("00000000000000000000000000000000"),	 -- 956	0
	 ("00000000000000000000000000000000"),	 -- 955	0
	 ("00000000000000000000000000000000"),	 -- 954	0
	 ("00000000000000000000000000000000"),	 -- 953	0
	 ("00000000000000000000000000000000"),	 -- 952	0
	 ("00000000000000000000000000000000"),	 -- 951	0
	 ("00000000000000000000000000000000"),	 -- 950	0
	 ("00000000000000000000000000000000"),	 -- 949	0
	 ("00000000000000000000000000000000"),	 -- 948	0
	 ("00000000000000000000000000000000"),	 -- 947	0
	 ("00000000000000000000000000000000"),	 -- 946	0
	 ("00000000000000000000000000000000"),	 -- 945	0
	 ("00000000000000000000000000000000"),	 -- 944	0
	 ("00000000000000000000000000000000"),	 -- 943	0
	 ("00000000000000000000000000000000"),	 -- 942	0
	 ("00000000000000000000000000000000"),	 -- 941	0
	 ("00000000000000000000000000000000"),	 -- 940	0
	 ("00000000000000000000000000000000"),	 -- 939	0
	 ("00000000000000000000000000000000"),	 -- 938	0
	 ("00000000000000000000000000000000"),	 -- 937	0
	 ("00000000000000000000000000000000"),	 -- 936	0
	 ("00000000000000000000000000000000"),	 -- 935	0
	 ("00000000000000000000000000000000"),	 -- 934	0
	 ("00000000000000000000000000000000"),	 -- 933	0
	 ("00000000000000000000000000000000"),	 -- 932	0
	 ("00000000000000000000000000000000"),	 -- 931	0
	 ("00000000000000000000000000000000"),	 -- 930	0
	 ("00000000000000000000000000000000"),	 -- 929	0
	 ("00000000000000000000000000000000"),	 -- 928	0
	 ("00000000000000000000000000000000"),	 -- 927	0
	 ("00000000000000000000000000000000"),	 -- 926	0
	 ("00000000000000000000000000000000"),	 -- 925	0
	 ("00000000000000000000000000000000"),	 -- 924	0
	 ("00000000000000000000000000000000"),	 -- 923	0
	 ("00000000000000000000000000000000"),	 -- 922	0
	 ("00000000000000000000000000000000"),	 -- 921	0
	 ("00000000000000000000000000000000"),	 -- 920	0
	 ("00000000000000000000000000000000"),	 -- 919	0
	 ("00000000000000000000000000000000"),	 -- 918	0
	 ("00000000000000000000000000000000"),	 -- 917	0
	 ("00000000000000000000000000000000"),	 -- 916	0
	 ("00000000000000000000000000000000"),	 -- 915	0
	 ("00000000000000000000000000000000"),	 -- 914	0
	 ("00000000000000000000000000000000"),	 -- 913	0
	 ("00000000000000000000000000000000"),	 -- 912	0
	 ("00000000000000000000000000000000"),	 -- 911	0
	 ("00000000000000000000000000000000"),	 -- 910	0
	 ("00000000000000000000000000000000"),	 -- 909	0
	 ("00000000000000000000000000000000"),	 -- 908	0
	 ("00000000000000000000000000000000"),	 -- 907	0
	 ("00000000000000000000000000000000"),	 -- 906	0
	 ("00000000000000000000000000000000"),	 -- 905	0
	 ("00000000000000000000000000000000"),	 -- 904	0
	 ("00000000000000000000000000000000"),	 -- 903	0
	 ("00000000000000000000000000000000"),	 -- 902	0
	 ("00000000000000000000000000000000"),	 -- 901	0
	 ("00000000000000000000000000000000"),	 -- 900	0
	 ("00000000000000000000000000000000"),	 -- 899	0
	 ("00000000000000000000000000000000"),	 -- 898	0
	 ("00000000000000000000000000000000"),	 -- 897	0
	 ("00000000000000000000000000000000"),	 -- 896	0
	 ("00000000000000000000000000000000"),	 -- 895	0
	 ("00000000000000000000000000000000"),	 -- 894	0
	 ("00000000000000000000000000000000"),	 -- 893	0
	 ("00000000000000000000000000000000"),	 -- 892	0
	 ("00000000000000000000000000000000"),	 -- 891	0
	 ("00000000000000000000000000000000"),	 -- 890	0
	 ("00000000000000000000000000000000"),	 -- 889	0
	 ("00000000000000000000000000000000"),	 -- 888	0
	 ("00000000000000000000000000000000"),	 -- 887	0
	 ("00000000000000000000000000000000"),	 -- 886	0
	 ("00000000000000000000000000000000"),	 -- 885	0
	 ("00000000000000000000000000000000"),	 -- 884	0
	 ("00000000000000000000000000000000"),	 -- 883	0
	 ("00000000000000000000000000000000"),	 -- 882	0
	 ("00000000000000000000000000000000"),	 -- 881	0
	 ("00000000000000000000000000000000"),	 -- 880	0
	 ("00000000000000000000000000000000"),	 -- 879	0
	 ("00000000000000000000000000000000"),	 -- 878	0
	 ("00000000000000000000000000000000"),	 -- 877	0
	 ("00000000000000000000000000000000"),	 -- 876	0
	 ("00000000000000000000000000000000"),	 -- 875	0
	 ("00000000000000000000000000000000"),	 -- 874	0
	 ("00000000000000000000000000000000"),	 -- 873	0
	 ("00000000000000000000000000000000"),	 -- 872	0
	 ("00000000000000000000000000000000"),	 -- 871	0
	 ("00000000000000000000000000000000"),	 -- 870	0
	 ("00000000000000000000000000000000"),	 -- 869	0
	 ("00000000000000000000000000000000"),	 -- 868	0
	 ("00000000000000000000000000000000"),	 -- 867	0
	 ("00000000000000000000000000000000"),	 -- 866	0
	 ("00000000000000000000000000000000"),	 -- 865	0
	 ("00000000000000000000000000000000"),	 -- 864	0
	 ("00000000000000000000000000000000"),	 -- 863	0
	 ("00000000000000000000000000000000"),	 -- 862	0
	 ("00000000000000000000000000000000"),	 -- 861	0
	 ("00000000000000000000000000000000"),	 -- 860	0
	 ("00000000000000000000000000000000"),	 -- 859	0
	 ("00000000000000000000000000000000"),	 -- 858	0
	 ("00000000000000000000000000000000"),	 -- 857	0
	 ("00000000000000000000000000000000"),	 -- 856	0
	 ("00000000000000000000000000000000"),	 -- 855	0
	 ("00000000000000000000000000000000"),	 -- 854	0
	 ("00000000000000000000000000000000"),	 -- 853	0
	 ("00000000000000000000000000000000"),	 -- 852	0
	 ("00000000000000000000000000000000"),	 -- 851	0
	 ("00000000000000000000000000000000"),	 -- 850	0
	 ("00000000000000000000000000000000"),	 -- 849	0
	 ("00000000000000000000000000000000"),	 -- 848	0
	 ("00000000000000000000000000000000"),	 -- 847	0
	 ("00000000000000000000000000000000"),	 -- 846	0
	 ("00000000000000000000000000000000"),	 -- 845	0
	 ("00000000000000000000000000000000"),	 -- 844	0
	 ("00000000000000000000000000000000"),	 -- 843	0
	 ("00000000000000000000000000000000"),	 -- 842	0
	 ("00000000000000000000000000000000"),	 -- 841	0
	 ("00000000000000000000000000000000"),	 -- 840	0
	 ("00000000000000000000000000000000"),	 -- 839	0
	 ("00000000000000000000000000000000"),	 -- 838	0
	 ("00000000000000000000000000000000"),	 -- 837	0
	 ("00000000000000000000000000000000"),	 -- 836	0
	 ("00000000000000000000000000000000"),	 -- 835	0
	 ("00000000000000000000000000000000"),	 -- 834	0
	 ("00000000000000000000000000000000"),	 -- 833	0
	 ("00000000000000000000000000000000"),	 -- 832	0
	 ("00000000000000000000000000000000"),	 -- 831	0
	 ("00000000000000000000000000000000"),	 -- 830	0
	 ("00000000000000000000000000000000"),	 -- 829	0
	 ("00000000000000000000000000000000"),	 -- 828	0
	 ("00000000000000000000000000000000"),	 -- 827	0
	 ("00000000000000000000000000000000"),	 -- 826	0
	 ("00000000000000000000000000000000"),	 -- 825	0
	 ("00000000000000000000000000000000"),	 -- 824	0
	 ("00000000000000000000000000000000"),	 -- 823	0
	 ("00000000000000000000000000000000"),	 -- 822	0
	 ("00000000000000000000000000000000"),	 -- 821	0
	 ("00000000000000000000000000000000"),	 -- 820	0
	 ("00000000000000000000000000000000"),	 -- 819	0
	 ("00000000000000000000000000000000"),	 -- 818	0
	 ("00000000000000000000000000000000"),	 -- 817	0
	 ("00000000000000000000000000000000"),	 -- 816	0
	 ("00000000000000000000000000000000"),	 -- 815	0
	 ("00000000000000000000000000000000"),	 -- 814	0
	 ("00000000000000000000000000000000"),	 -- 813	0
	 ("00000000000000000000000000000000"),	 -- 812	0
	 ("00000000000000000000000000000000"),	 -- 811	0
	 ("00000000000000000000000000000000"),	 -- 810	0
	 ("00000000000000000000000000000000"),	 -- 809	0
	 ("00000000000000000000000000000000"),	 -- 808	0
	 ("00000000000000000000000000000000"),	 -- 807	0
	 ("00000000000000000000000000000000"),	 -- 806	0
	 ("00000000000000000000000000000000"),	 -- 805	0
	 ("00000000000000000000000000000000"),	 -- 804	0
	 ("00000000000000000000000000000000"),	 -- 803	0
	 ("00000000000000000000000000000000"),	 -- 802	0
	 ("00000000000000000000000000000000"),	 -- 801	0
	 ("00000000000000000000000000000000"),	 -- 800	0
	 ("00000000000000000000000000000000"),	 -- 799	0
	 ("00000000000000000000000000000000"),	 -- 798	0
	 ("00000000000000000000000000000000"),	 -- 797	0
	 ("00000000000000000000000000000000"),	 -- 796	0
	 ("00000000000000000000000000000000"),	 -- 795	0
	 ("00000000000000000000000000000000"),	 -- 794	0
	 ("00000000000000000000000000000000"),	 -- 793	0
	 ("00000000000000000000000000000000"),	 -- 792	0
	 ("00000000000000000000000000000000"),	 -- 791	0
	 ("00000000000000000000000000000000"),	 -- 790	0
	 ("00000000000000000000000000000000"),	 -- 789	0
	 ("00000000000000000000000000000000"),	 -- 788	0
	 ("00000000000000000000000000000000"),	 -- 787	0
	 ("00000000000000000000000000000000"),	 -- 786	0
	 ("00000000000000000000000000000000"),	 -- 785	0
	 ("00000000000000000000000000000000"),	 -- 784	0
	 ("00000000000000000000000000000000"),	 -- 783	0
	 ("00000000000000000000000000000000"),	 -- 782	0
	 ("00000000000000000000000000000000"),	 -- 781	0
	 ("00000000000000000000000000000000"),	 -- 780	0
	 ("00000000000000000000000000000000"),	 -- 779	0
	 ("00000000000000000000000000000000"),	 -- 778	0
	 ("00000000000000000000000000000000"),	 -- 777	0
	 ("00000000000000000000000000000000"),	 -- 776	0
	 ("00000000000000000000000000000000"),	 -- 775	0
	 ("00000000000000000000000000000000"),	 -- 774	0
	 ("00000000000000000000000000000000"),	 -- 773	0
	 ("00000000000000000000000000000000"),	 -- 772	0
	 ("00000000000000000000000000000000"),	 -- 771	0
	 ("00000000000000000000000000000000"),	 -- 770	0
	 ("00000000000000000000000000000000"),	 -- 769	0
	 ("00000000000000000000000000000000"),	 -- 768	0
	 ("00000000000000000000000000000000"),	 -- 767	0
	 ("00000000000000000000000000000000"),	 -- 766	0
	 ("00000000000000000000000000000000"),	 -- 765	0
	 ("00000000000000000000000000000000"),	 -- 764	0
	 ("00000000000000000000000000000000"),	 -- 763	0
	 ("00000000000000000000000000000000"),	 -- 762	0
	 ("00000000000000000000000000000000"),	 -- 761	0
	 ("00000000000000000000000000000000"),	 -- 760	0
	 ("00000000000000000000000000000000"),	 -- 759	0
	 ("00000000000000000000000000000000"),	 -- 758	0
	 ("00000000000000000000000000000000"),	 -- 757	0
	 ("00000000000000000000000000000000"),	 -- 756	0
	 ("00000000000000000000000000000000"),	 -- 755	0
	 ("00000000000000000000000000000000"),	 -- 754	0
	 ("00000000000000000000000000000000"),	 -- 753	0
	 ("00000000000000000000000000000000"),	 -- 752	0
	 ("00000000000000000000000000000000"),	 -- 751	0
	 ("00000000000000000000000000000000"),	 -- 750	0
	 ("00000000000000000000000000000000"),	 -- 749	0
	 ("00000000000000000000000000000000"),	 -- 748	0
	 ("00000000000000000000000000000000"),	 -- 747	0
	 ("00000000000000000000000000000000"),	 -- 746	0
	 ("00000000000000000000000000000000"),	 -- 745	0
	 ("00000000000000000000000000000000"),	 -- 744	0
	 ("00000000000000000000000000000000"),	 -- 743	0
	 ("00000000000000000000000000000000"),	 -- 742	0
	 ("00000000000000000000000000000000"),	 -- 741	0
	 ("00000000000000000000000000000000"),	 -- 740	0
	 ("00000000000000000000000000000000"),	 -- 739	0
	 ("00000000000000000000000000000000"),	 -- 738	0
	 ("00000000000000000000000000000000"),	 -- 737	0
	 ("00000000000000000000000000000000"),	 -- 736	0
	 ("00000000000000000000000000000000"),	 -- 735	0
	 ("00000000000000000000000000000000"),	 -- 734	0
	 ("00000000000000000000000000000000"),	 -- 733	0
	 ("00000000000000000000000000000000"),	 -- 732	0
	 ("00000000000000000000000000000000"),	 -- 731	0
	 ("00000000000000000000000000000000"),	 -- 730	0
	 ("00000000000000000000000000000000"),	 -- 729	0
	 ("00000000000000000000000000000000"),	 -- 728	0
	 ("00000000000000000000000000000000"),	 -- 727	0
	 ("00000000000000000000000000000000"),	 -- 726	0
	 ("00000000000000000000000000000000"),	 -- 725	0
	 ("00000000000000000000000000000000"),	 -- 724	0
	 ("00000000000000000000000000000000"),	 -- 723	0
	 ("00000000000000000000000000000000"),	 -- 722	0
	 ("00000000000000000000000000000000"),	 -- 721	0
	 ("00000000000000000000000000000000"),	 -- 720	0
	 ("00000000000000000000000000000000"),	 -- 719	0
	 ("00000000000000000000000000000000"),	 -- 718	0
	 ("00000000000000000000000000000000"),	 -- 717	0
	 ("00000000000000000000000000000000"),	 -- 716	0
	 ("00000000000000000000000000000000"),	 -- 715	0
	 ("00000000000000000000000000000000"),	 -- 714	0
	 ("00000000000000000000000000000000"),	 -- 713	0
	 ("00000000000000000000000000000000"),	 -- 712	0
	 ("00000000000000000000000000000000"),	 -- 711	0
	 ("00000000000000000000000000000000"),	 -- 710	0
	 ("00000000000000000000000000000000"),	 -- 709	0
	 ("00000000000000000000000000000000"),	 -- 708	0
	 ("00000000000000000000000000000000"),	 -- 707	0
	 ("00000000000000000000000000000000"),	 -- 706	0
	 ("00000000000000000000000000000000"),	 -- 705	0
	 ("00000000000000000000000000000000"),	 -- 704	0
	 ("00000000000000000000000000000000"),	 -- 703	0
	 ("00000000000000000000000000000000"),	 -- 702	0
	 ("00000000000000000000000000000000"),	 -- 701	0
	 ("00000000000000000000000000000000"),	 -- 700	0
	 ("00000000000000000000000000000000"),	 -- 699	0
	 ("00000000000000000000000000000000"),	 -- 698	0
	 ("00000000000000000000000000000000"),	 -- 697	0
	 ("00000000000000000000000000000000"),	 -- 696	0
	 ("00000000000000000000000000000000"),	 -- 695	0
	 ("00000000000000000000000000000000"),	 -- 694	0
	 ("00000000000000000000000000000000"),	 -- 693	0
	 ("00000000000000000000000000000000"),	 -- 692	0
	 ("00000000000000000000000000000000"),	 -- 691	0
	 ("00000000000000000000000000000000"),	 -- 690	0
	 ("00000000000000000000000000000000"),	 -- 689	0
	 ("00000000000000000000000000000000"),	 -- 688	0
	 ("00000000000000000000000000000000"),	 -- 687	0
	 ("00000000000000000000000000000000"),	 -- 686	0
	 ("00000000000000000000000000000000"),	 -- 685	0
	 ("00000000000000000000000000000000"),	 -- 684	0
	 ("00000000000000000000000000000000"),	 -- 683	0
	 ("00000000000000000000000000000000"),	 -- 682	0
	 ("00000000000000000000000000000000"),	 -- 681	0
	 ("00000000000000000000000000000000"),	 -- 680	0
	 ("00000000000000000000000000000000"),	 -- 679	0
	 ("00000000000000000000000000000000"),	 -- 678	0
	 ("00000000000000000000000000000000"),	 -- 677	0
	 ("00000000000000000000000000000000"),	 -- 676	0
	 ("00000000000000000000000000000000"),	 -- 675	0
	 ("00000000000000000000000000000000"),	 -- 674	0
	 ("00000000000000000000000000000000"),	 -- 673	0
	 ("00000000000000000000000000000000"),	 -- 672	0
	 ("00000000000000000000000000000000"),	 -- 671	0
	 ("00000000000000000000000000000000"),	 -- 670	0
	 ("00000000000000000000000000000000"),	 -- 669	0
	 ("00000000000000000000000000000000"),	 -- 668	0
	 ("00000000000000000000000000000000"),	 -- 667	0
	 ("00000000000000000000000000000000"),	 -- 666	0
	 ("00000000000000000000000000000000"),	 -- 665	0
	 ("00000000000000000000000000000000"),	 -- 664	0
	 ("00000000000000000000000000000000"),	 -- 663	0
	 ("00000000000000000000000000000000"),	 -- 662	0
	 ("00000000000000000000000000000000"),	 -- 661	0
	 ("00000000000000000000000000000000"),	 -- 660	0
	 ("00000000000000000000000000000000"),	 -- 659	0
	 ("00000000000000000000000000000000"),	 -- 658	0
	 ("00000000000000000000000000000000"),	 -- 657	0
	 ("00000000000000000000000000000000"),	 -- 656	0
	 ("00000000000000000000000000000000"),	 -- 655	0
	 ("00000000000000000000000000000000"),	 -- 654	0
	 ("00000000000000000000000000000000"),	 -- 653	0
	 ("00000000000000000000000000000000"),	 -- 652	0
	 ("00000000000000000000000000000000"),	 -- 651	0
	 ("00000000000000000000000000000000"),	 -- 650	0
	 ("00000000000000000000000000000000"),	 -- 649	0
	 ("00000000000000000000000000000000"),	 -- 648	0
	 ("00000000000000000000000000000000"),	 -- 647	0
	 ("00000000000000000000000000000000"),	 -- 646	0
	 ("00000000000000000000000000000000"),	 -- 645	0
	 ("00000000000000000000000000000000"),	 -- 644	0
	 ("00000000000000000000000000000000"),	 -- 643	0
	 ("00000000000000000000000000000000"),	 -- 642	0
	 ("00000000000000000000000000000000"),	 -- 641	0
	 ("00000000000000000000000000000000"),	 -- 640	0
	 ("00000000000000000000000000000000"),	 -- 639	0
	 ("00000000000000000000000000000000"),	 -- 638	0
	 ("00000000000000000000000000000000"),	 -- 637	0
	 ("00000000000000000000000000000000"),	 -- 636	0
	 ("00000000000000000000000000000000"),	 -- 635	0
	 ("00000000000000000000000000000000"),	 -- 634	0
	 ("00000000000000000000000000000000"),	 -- 633	0
	 ("00000000000000000000000000000000"),	 -- 632	0
	 ("00000000000000000000000000000000"),	 -- 631	0
	 ("00000000000000000000000000000000"),	 -- 630	0
	 ("00000000000000000000000000000000"),	 -- 629	0
	 ("00000000000000000000000000000000"),	 -- 628	0
	 ("00000000000000000000000000000000"),	 -- 627	0
	 ("00000000000000000000000000000000"),	 -- 626	0
	 ("00000000000000000000000000000000"),	 -- 625	0
	 ("00000000000000000000000000000000"),	 -- 624	0
	 ("00000000000000000000000000000000"),	 -- 623	0
	 ("00000000000000000000000000000000"),	 -- 622	0
	 ("00000000000000000000000000000000"),	 -- 621	0
	 ("00000000000000000000000000000000"),	 -- 620	0
	 ("00000000000000000000000000000000"),	 -- 619	0
	 ("00000000000000000000000000000000"),	 -- 618	0
	 ("00000000000000000000000000000000"),	 -- 617	0
	 ("00000000000000000000000000000000"),	 -- 616	0
	 ("00000000000000000000000000000000"),	 -- 615	0
	 ("00000000000000000000000000000000"),	 -- 614	0
	 ("00000000000000000000000000000000"),	 -- 613	0
	 ("00000000000000000000000000000000"),	 -- 612	0
	 ("00000000000000000000000000000000"),	 -- 611	0
	 ("00000000000000000000000000000000"),	 -- 610	0
	 ("00000000000000000000000000000000"),	 -- 609	0
	 ("00000000000000000000000000000000"),	 -- 608	0
	 ("00000000000000000000000000000000"),	 -- 607	0
	 ("00000000000000000000000000000000"),	 -- 606	0
	 ("00000000000000000000000000000000"),	 -- 605	0
	 ("00000000000000000000000000000000"),	 -- 604	0
	 ("00000000000000000000000000000000"),	 -- 603	0
	 ("00000000000000000000000000000000"),	 -- 602	0
	 ("00000000000000000000000000000000"),	 -- 601	0
	 ("00000000000000000000000000000000"),	 -- 600	0
	 ("00000000000000000000000000000000"),	 -- 599	0
	 ("00000000000000000000000000000000"),	 -- 598	0
	 ("00000000000000000000000000000000"),	 -- 597	0
	 ("00000000000000000000000000000000"),	 -- 596	0
	 ("00000000000000000000000000000000"),	 -- 595	0
	 ("00000000000000000000000000000000"),	 -- 594	0
	 ("00000000000000000000000000000000"),	 -- 593	0
	 ("00000000000000000000000000000000"),	 -- 592	0
	 ("00000000000000000000000000000000"),	 -- 591	0
	 ("00000000000000000000000000000000"),	 -- 590	0
	 ("00000000000000000000000000000000"),	 -- 589	0
	 ("00000000000000000000000000000000"),	 -- 588	0
	 ("00000000000000000000000000000000"),	 -- 587	0
	 ("00000000000000000000000000000000"),	 -- 586	0
	 ("00000000000000000000000000000000"),	 -- 585	0
	 ("00000000000000000000000000000000"),	 -- 584	0
	 ("00000000000000000000000000000000"),	 -- 583	0
	 ("00000000000000000000000000000000"),	 -- 582	0
	 ("00000000000000000000000000000000"),	 -- 581	0
	 ("00000000000000000000000000000000"),	 -- 580	0
	 ("00000000000000000000000000000000"),	 -- 579	0
	 ("00000000000000000000000000000000"),	 -- 578	0
	 ("00000000000000000000000000000000"),	 -- 577	0
	 ("00000000000000000000000000000000"),	 -- 576	0
	 ("00000000000000000000000000000000"),	 -- 575	0
	 ("00000000000000000000000000000000"),	 -- 574	0
	 ("00000000000000000000000000000000"),	 -- 573	0
	 ("00000000000000000000000000000000"),	 -- 572	0
	 ("00000000000000000000000000000000"),	 -- 571	0
	 ("00000000000000000000000000000000"),	 -- 570	0
	 ("00000000000000000000000000000000"),	 -- 569	0
	 ("00000000000000000000000000000000"),	 -- 568	0
	 ("00000000000000000000000000000000"),	 -- 567	0
	 ("00000000000000000000000000000000"),	 -- 566	0
	 ("00000000000000000000000000000000"),	 -- 565	0
	 ("00000000000000000000000000000000"),	 -- 564	0
	 ("00000000000000000000000000000000"),	 -- 563	0
	 ("00000000000000000000000000000000"),	 -- 562	0
	 ("00000000000000000000000000000000"),	 -- 561	0
	 ("00000000000000000000000000000000"),	 -- 560	0
	 ("00000000000000000000000000000000"),	 -- 559	0
	 ("00000000000000000000000000000000"),	 -- 558	0
	 ("00000000000000000000000000000000"),	 -- 557	0
	 ("00000000000000000000000000000000"),	 -- 556	0
	 ("00000000000000000000000000000000"),	 -- 555	0
	 ("00000000000000000000000000000000"),	 -- 554	0
	 ("00000000000000000000000000000000"),	 -- 553	0
	 ("00000000000000000000000000000000"),	 -- 552	0
	 ("00000000000000000000000000000000"),	 -- 551	0
	 ("00000000000000000000000000000000"),	 -- 550	0
	 ("00000000000000000000000000000000"),	 -- 549	0
	 ("00000000000000000000000000000000"),	 -- 548	0
	 ("00000000000000000000000000000000"),	 -- 547	0
	 ("00000000000000000000000000000000"),	 -- 546	0
	 ("00000000000000000000000000000000"),	 -- 545	0
	 ("00000000000000000000000000000000"),	 -- 544	0
	 ("00000000000000000000000000000000"),	 -- 543	0
	 ("00000000000000000000000000000000"),	 -- 542	0
	 ("00000000000000000000000000000000"),	 -- 541	0
	 ("00000000000000000000000000000000"),	 -- 540	0
	 ("00000000000000000000000000000000"),	 -- 539	0
	 ("00000000000000000000000000000000"),	 -- 538	0
	 ("00000000000000000000000000000000"),	 -- 537	0
	 ("00000000000000000000000000000000"),	 -- 536	0
	 ("00000000000000000000000000000000"),	 -- 535	0
	 ("00000000000000000000000000000000"),	 -- 534	0
	 ("00000000000000000000000000000000"),	 -- 533	0
	 ("00000000000000000000000000000000"),	 -- 532	0
	 ("00000000000000000000000000000000"),	 -- 531	0
	 ("00000000000000000000000000000000"),	 -- 530	0
	 ("00000000000000000000000000000000"),	 -- 529	0
	 ("00000000000000000000000000000000"),	 -- 528	0
	 ("00000000000000000000000000000000"),	 -- 527	0
	 ("00000000000000000000000000000000"),	 -- 526	0
	 ("00000000000000000000000000000000"),	 -- 525	0
	 ("00000000000000000000000000000000"),	 -- 524	0
	 ("00000000000000000000000000000000"),	 -- 523	0
	 ("00000000000000000000000000000000"),	 -- 522	0
	 ("00000000000000000000000000000000"),	 -- 521	0
	 ("00000000000000000000000000000000"),	 -- 520	0
	 ("00000000000000000000000000000000"),	 -- 519	0
	 ("00000000000000000000000000000000"),	 -- 518	0
	 ("00000000000000000000000000000000"),	 -- 517	0
	 ("00000000000000000000000000000000"),	 -- 516	0
	 ("00000000000000000000000000000000"),	 -- 515	0
	 ("00000000000000000000000000000000"),	 -- 514	0
	 ("00000000000000000000000000000000"),	 -- 513	0
	 ("00000000000000000000000000000000"),	 -- 512	0
	 ("00000000000000000000000000000000"),	 -- 511	0
	 ("00000000000000000000000000000000"),	 -- 510	0
	 ("00000000000000000000000000000000"),	 -- 509	0
	 ("00000000000000000000000000000000"),	 -- 508	0
	 ("00000000000000000000000000000000"),	 -- 507	0
	 ("00000000000000000000000000000000"),	 -- 506	0
	 ("00000000000000000000000000000000"),	 -- 505	0
	 ("00000000000000000000000000000000"),	 -- 504	0
	 ("00000000000000000000000000000000"),	 -- 503	0
	 ("00000000000000000000000000000000"),	 -- 502	0
	 ("00000000000000000000000000000000"),	 -- 501	0
	 ("00000000000000000000000000000000"),	 -- 500	0
	 ("00000000000000000000000000000000"),	 -- 499	0
	 ("00000000000000000000000000000000"),	 -- 498	0
	 ("00000000000000000000000000000000"),	 -- 497	0
	 ("00000000000000000000000000000000"),	 -- 496	0
	 ("00000000000000000000000000000000"),	 -- 495	0
	 ("00000000000000000000000000000000"),	 -- 494	0
	 ("00000000000000000000000000000000"),	 -- 493	0
	 ("00000000000000000000000000000000"),	 -- 492	0
	 ("00000000000000000000000000000000"),	 -- 491	0
	 ("00000000000000000000000000000000"),	 -- 490	0
	 ("00000000000000000000000000000000"),	 -- 489	0
	 ("00000000000000000000000000000000"),	 -- 488	0
	 ("00000000000000000000000000000000"),	 -- 487	0
	 ("00000000000000000000000000000000"),	 -- 486	0
	 ("00000000000000000000000000000000"),	 -- 485	0
	 ("00000000000000000000000000000000"),	 -- 484	0
	 ("00000000000000000000000000000000"),	 -- 483	0
	 ("00000000000000000000000000000000"),	 -- 482	0
	 ("00000000000000000000000000000000"),	 -- 481	0
	 ("00000000000000000000000000000000"),	 -- 480	0
	 ("00000000000000000000000000000000"),	 -- 479	0
	 ("00000000000000000000000000000000"),	 -- 478	0
	 ("00000000000000000000000000000000"),	 -- 477	0
	 ("00000000000000000000000000000000"),	 -- 476	0
	 ("00000000000000000000000000000000"),	 -- 475	0
	 ("00000000000000000000000000000000"),	 -- 474	0
	 ("00000000000000000000000000000000"),	 -- 473	0
	 ("00000000000000000000000000000000"),	 -- 472	0
	 ("00000000000000000000000000000000"),	 -- 471	0
	 ("00000000000000000000000000000000"),	 -- 470	0
	 ("00000000000000000000000000000000"),	 -- 469	0
	 ("00000000000000000000000000000000"),	 -- 468	0
	 ("00000000000000000000000000000000"),	 -- 467	0
	 ("00000000000000000000000000000000"),	 -- 466	0
	 ("00000000000000000000000000000000"),	 -- 465	0
	 ("00000000000000000000000000000000"),	 -- 464	0
	 ("00000000000000000000000000000000"),	 -- 463	0
	 ("00000000000000000000000000000000"),	 -- 462	0
	 ("00000000000000000000000000000000"),	 -- 461	0
	 ("00000000000000000000000000000000"),	 -- 460	0
	 ("00000000000000000000000000000000"),	 -- 459	0
	 ("00000000000000000000000000000000"),	 -- 458	0
	 ("00000000000000000000000000000000"),	 -- 457	0
	 ("00000000000000000000000000000000"),	 -- 456	0
	 ("00000000000000000000000000000000"),	 -- 455	0
	 ("00000000000000000000000000000000"),	 -- 454	0
	 ("00000000000000000000000000000000"),	 -- 453	0
	 ("00000000000000000000000000000000"),	 -- 452	0
	 ("00000000000000000000000000000000"),	 -- 451	0
	 ("00000000000000000000000000000000"),	 -- 450	0
	 ("00000000000000000000000000000000"),	 -- 449	0
	 ("00000000000000000000000000000000"),	 -- 448	0
	 ("00000000000000000000000000000000"),	 -- 447	0
	 ("00000000000000000000000000000000"),	 -- 446	0
	 ("00000000000000000000000000000000"),	 -- 445	0
	 ("00000000000000000000000000000000"),	 -- 444	0
	 ("00000000000000000000000000000000"),	 -- 443	0
	 ("00000000000000000000000000000000"),	 -- 442	0
	 ("00000000000000000000000000000000"),	 -- 441	0
	 ("00000000000000000000000000000000"),	 -- 440	0
	 ("00000000000000000000000000000000"),	 -- 439	0
	 ("00000000000000000000000000000000"),	 -- 438	0
	 ("00000000000000000000000000000000"),	 -- 437	0
	 ("00000000000000000000000000000000"),	 -- 436	0
	 ("00000000000000000000000000000000"),	 -- 435	0
	 ("00000000000000000000000000000000"),	 -- 434	0
	 ("00000000000000000000000000000000"),	 -- 433	0
	 ("00000000000000000000000000000000"),	 -- 432	0
	 ("00000000000000000000000000000000"),	 -- 431	0
	 ("00000000000000000000000000000000"),	 -- 430	0
	 ("00000000000000000000000000000000"),	 -- 429	0
	 ("00000000000000000000000000000000"),	 -- 428	0
	 ("00000000000000000000000000000000"),	 -- 427	0
	 ("00000000000000000000000000000000"),	 -- 426	0
	 ("00000000000000000000000000000000"),	 -- 425	0
	 ("00000000000000000000000000000000"),	 -- 424	0
	 ("00000000000000000000000000000000"),	 -- 423	0
	 ("00000000000000000000000000000000"),	 -- 422	0
	 ("00000000000000000000000000000000"),	 -- 421	0
	 ("00000000000000000000000000000000"),	 -- 420	0
	 ("00000000000000000000000000000000"),	 -- 419	0
	 ("00000000000000000000000000000000"),	 -- 418	0
	 ("00000000000000000000000000000000"),	 -- 417	0
	 ("00000000000000000000000000000000"),	 -- 416	0
	 ("00000000000000000000000000000000"),	 -- 415	0
	 ("00000000000000000000000000000000"),	 -- 414	0
	 ("00000000000000000000000000000000"),	 -- 413	0
	 ("00000000000000000000000000000000"),	 -- 412	0
	 ("00000000000000000000000000000000"),	 -- 411	0
	 ("00000000000000000000000000000000"),	 -- 410	0
	 ("00000000000000000000000000000000"),	 -- 409	0
	 ("00000000000000000000000000000000"),	 -- 408	0
	 ("00000000000000000000000000000000"),	 -- 407	0
	 ("00000000000000000000000000000000"),	 -- 406	0
	 ("00000000000000000000000000000000"),	 -- 405	0
	 ("00000000000000000000000000000000"),	 -- 404	0
	 ("00000000000000000000000000000000"),	 -- 403	0
	 ("00000000000000000000000000000000"),	 -- 402	0
	 ("00000000000000000000000000000000"),	 -- 401	0
	 ("00000000000000000000000000000000"),	 -- 400	0
	 ("00000000000000000000000000000000"),	 -- 399	0
	 ("00000000000000000000000000000000"),	 -- 398	0
	 ("00000000000000000000000000000000"),	 -- 397	0
	 ("00000000000000000000000000000000"),	 -- 396	0
	 ("00000000000000000000000000000000"),	 -- 395	0
	 ("00000000000000000000000000000000"),	 -- 394	0
	 ("00000000000000000000000000000000"),	 -- 393	0
	 ("00000000000000000000000000000000"),	 -- 392	0
	 ("00000000000000000000000000000000"),	 -- 391	0
	 ("00000000000000000000000000000000"),	 -- 390	0
	 ("00000000000000000000000000000000"),	 -- 389	0
	 ("00000000000000000000000000000000"),	 -- 388	0
	 ("00000000000000000000000000000000"),	 -- 387	0
	 ("00000000000000000000000000000000"),	 -- 386	0
	 ("00000000000000000000000000000000"),	 -- 385	0
	 ("00000000000000000000000000000000"),	 -- 384	0
	 ("00000000000000000000000000000000"),	 -- 383	0
	 ("00000000000000000000000000000000"),	 -- 382	0
	 ("00000000000000000000000000000000"),	 -- 381	0
	 ("00000000000000000000000000000000"),	 -- 380	0
	 ("00000000000000000000000000000000"),	 -- 379	0
	 ("00000000000000000000000000000000"),	 -- 378	0
	 ("00000000000000000000000000000000"),	 -- 377	0
	 ("00000000000000000000000000000000"),	 -- 376	0
	 ("00000000000000000000000000000000"),	 -- 375	0
	 ("00000000000000000000000000000000"),	 -- 374	0
	 ("00000000000000000000000000000000"),	 -- 373	0
	 ("00000000000000000000000000000000"),	 -- 372	0
	 ("00000000000000000000000000000000"),	 -- 371	0
	 ("00000000000000000000000000000000"),	 -- 370	0
	 ("00000000000000000000000000000000"),	 -- 369	0
	 ("00000000000000000000000000000000"),	 -- 368	0
	 ("00000000000000000000000000000000"),	 -- 367	0
	 ("00000000000000000000000000000000"),	 -- 366	0
	 ("00000000000000000000000000000000"),	 -- 365	0
	 ("00000000000000000000000000000000"),	 -- 364	0
	 ("00000000000000000000000000000000"),	 -- 363	0
	 ("00000000000000000000000000000000"),	 -- 362	0
	 ("00000000000000000000000000000000"),	 -- 361	0
	 ("00000000000000000000000000000000"),	 -- 360	0
	 ("00000000000000000000000000000000"),	 -- 359	0
	 ("00000000000000000000000000000000"),	 -- 358	0
	 ("00000000000000000000000000000000"),	 -- 357	0
	 ("00000000000000000000000000000000"),	 -- 356	0
	 ("00000000000000000000000000000000"),	 -- 355	0
	 ("00000000000000000000000000000000"),	 -- 354	0
	 ("00000000000000000000000000000000"),	 -- 353	0
	 ("00000000000000000000000000000000"),	 -- 352	0
	 ("00000000000000000000000000000000"),	 -- 351	0
	 ("00000000000000000000000000000000"),	 -- 350	0
	 ("00000000000000000000000000000000"),	 -- 349	0
	 ("00000000000000000000000000000000"),	 -- 348	0
	 ("00000000000000000000000000000000"),	 -- 347	0
	 ("00000000000000000000000000000000"),	 -- 346	0
	 ("00000000000000000000000000000000"),	 -- 345	0
	 ("00000000000000000000000000000000"),	 -- 344	0
	 ("00000000000000000000000000000000"),	 -- 343	0
	 ("00000000000000000000000000000000"),	 -- 342	0
	 ("00000000000000000000000000000000"),	 -- 341	0
	 ("00000000000000000000000000000000"),	 -- 340	0
	 ("00000000000000000000000000000000"),	 -- 339	0
	 ("00000000000000000000000000000000"),	 -- 338	0
	 ("00000000000000000000000000000000"),	 -- 337	0
	 ("00000000000000000000000000000000"),	 -- 336	0
	 ("00000000000000000000000000000000"),	 -- 335	0
	 ("00000000000000000000000000000000"),	 -- 334	0
	 ("00000000000000000000000000000000"),	 -- 333	0
	 ("00000000000000000000000000000000"),	 -- 332	0
	 ("00000000000000000000000000000000"),	 -- 331	0
	 ("00000000000000000000000000000000"),	 -- 330	0
	 ("00000000000000000000000000000000"),	 -- 329	0
	 ("00000000000000000000000000000000"),	 -- 328	0
	 ("00000000000000000000000000000000"),	 -- 327	0
	 ("00000000000000000000000000000000"),	 -- 326	0
	 ("00000000000000000000000000000000"),	 -- 325	0
	 ("00000000000000000000000000000000"),	 -- 324	0
	 ("00000000000000000000000000000000"),	 -- 323	0
	 ("00000000000000000000000000000000"),	 -- 322	0
	 ("00000000000000000000000000000000"),	 -- 321	0
	 ("00000000000000000000000000000000"),	 -- 320	0
	 ("00000000000000000000000000000000"),	 -- 319	0
	 ("00000000000000000000000000000000"),	 -- 318	0
	 ("00000000000000000000000000000000"),	 -- 317	0
	 ("00000000000000000000000000000000"),	 -- 316	0
	 ("00000000000000000000000000000000"),	 -- 315	0
	 ("00000000000000000000000000000000"),	 -- 314	0
	 ("00000000000000000000000000000000"),	 -- 313	0
	 ("00000000000000000000000000000000"),	 -- 312	0
	 ("00000000000000000000000000000000"),	 -- 311	0
	 ("00000000000000000000000000000000"),	 -- 310	0
	 ("00000000000000000000000000000000"),	 -- 309	0
	 ("00000000000000000000000000000000"),	 -- 308	0
	 ("00000000000000000000000000000000"),	 -- 307	0
	 ("00000000000000000000000000000000"),	 -- 306	0
	 ("00000000000000000000000000000000"),	 -- 305	0
	 ("00000000000000000000000000000000"),	 -- 304	0
	 ("00000000000000000000000000000000"),	 -- 303	0
	 ("00000000000000000000000000000000"),	 -- 302	0
	 ("00000000000000000000000000000000"),	 -- 301	0
	 ("00000000000000000000000000000000"),	 -- 300	0
	 ("00000000000000000000000000000000"),	 -- 299	0
	 ("00000000000000000000000000000000"),	 -- 298	0
	 ("00000000000000000000000000000000"),	 -- 297	0
	 ("00000000000000000000000000000000"),	 -- 296	0
	 ("00000000000000000000000000000000"),	 -- 295	0
	 ("00000000000000000000000000000000"),	 -- 294	0
	 ("00000000000000000000000000000000"),	 -- 293	0
	 ("00000000000000000000000000000000"),	 -- 292	0
	 ("00000000000000000000000000000000"),	 -- 291	0
	 ("00000000000000000000000000000000"),	 -- 290	0
	 ("00000000000000000000000000000000"),	 -- 289	0
	 ("00000000000000000000000000000000"),	 -- 288	0
	 ("00000000000000000000000000000000"),	 -- 287	0
	 ("00000000000000000000000000000000"),	 -- 286	0
	 ("00000000000000000000000000000000"),	 -- 285	0
	 ("00000000000000000000000000000000"),	 -- 284	0
	 ("00000000000000000000000000000000"),	 -- 283	0
	 ("00000000000000000000000000000000"),	 -- 282	0
	 ("00000000000000000000000000000000"),	 -- 281	0
	 ("00000000000000000000000000000000"),	 -- 280	0
	 ("00000000000000000000000000000000"),	 -- 279	0
	 ("00000000000000000000000000000000"),	 -- 278	0
	 ("00000000000000000000000000000000"),	 -- 277	0
	 ("00000000000000000000000000000000"),	 -- 276	0
	 ("00000000000000000000000000000000"),	 -- 275	0
	 ("00000000000000000000000000000000"),	 -- 274	0
	 ("00000000000000000000000000000000"),	 -- 273	0
	 ("00000000000000000000000000000000"),	 -- 272	0
	 ("00000000000000000000000000000000"),	 -- 271	0
	 ("00000000000000000000000000000000"),	 -- 270	0
	 ("00000000000000000000000000000000"),	 -- 269	0
	 ("00000000000000000000000000000000"),	 -- 268	0
	 ("00000000000000000000000000000000"),	 -- 267	0
	 ("00000000000000000000000000000000"),	 -- 266	0
	 ("00000000000000000000000000000000"),	 -- 265	0
	 ("00000000000000000000000000000000"),	 -- 264	0
	 ("00000000000000000000000000000000"),	 -- 263	0
	 ("00000000000000000000000000000000"),	 -- 262	0
	 ("00000000000000000000000000000000"),	 -- 261	0
	 ("00000000000000000000000000000000"),	 -- 260	0
	 ("00000000000000000000000000000000"),	 -- 259	0
	 ("00000000000000000000000000000000"),	 -- 258	0
	 ("00000000000000000000000000000000"),	 -- 257	0
	 ("00000000000000000000000000000000"),	 -- 256	0
	 ("00000000000000000000000000000000"),	 -- 255	0
	 ("00000000000000000000000000000000"),	 -- 254	0
	 ("00000000000000000000000000000000"),	 -- 253	0
	 ("00000000000000000000000000000000"),	 -- 252	0
	 ("00000000000000000000000000000000"),	 -- 251	0
	 ("00000000000000000000000000000000"),	 -- 250	0
	 ("00000000000000000000000000000000"),	 -- 249	0
	 ("00000000000000000000000000000000"),	 -- 248	0
	 ("00000000000000000000000000000000"),	 -- 247	0
	 ("00000000000000000000000000000000"),	 -- 246	0
	 ("00000000000000000000000000000000"),	 -- 245	0
	 ("00000000000000000000000000000000"),	 -- 244	0
	 ("00000000000000000000000000000000"),	 -- 243	0
	 ("00000000000000000000000000000000"),	 -- 242	0
	 ("00000000000000000000000000000000"),	 -- 241	0
	 ("00000000000000000000000000000000"),	 -- 240	0
	 ("00000000000000000000000000000000"),	 -- 239	0
	 ("00000000000000000000000000000000"),	 -- 238	0
	 ("00000000000000000000000000000000"),	 -- 237	0
	 ("00000000000000000000000000000000"),	 -- 236	0
	 ("00000000000000000000000000000000"),	 -- 235	0
	 ("00000000000000000000000000000000"),	 -- 234	0
	 ("00000000000000000000000000000000"),	 -- 233	0
	 ("00000000000000000000000000000000"),	 -- 232	0
	 ("00000000000000000000000000000000"),	 -- 231	0
	 ("00000000000000000000000000000000"),	 -- 230	0
	 ("00000000000000000000000000000000"),	 -- 229	0
	 ("00000000000000000000000000000000"),	 -- 228	0
	 ("00000000000000000000000000000000"),	 -- 227	0
	 ("00000000000000000000000000000000"),	 -- 226	0
	 ("00000000000000000000000000000000"),	 -- 225	0
	 ("00000000000000000000000000000000"),	 -- 224	0
	 ("00000000000000000000000000000000"),	 -- 223	0
	 ("00000000000000000000000000000000"),	 -- 222	0
	 ("00000000000000000000000000000000"),	 -- 221	0
	 ("00000000000000000000000000000000"),	 -- 220	0
	 ("00000000000000000000000000000000"),	 -- 219	0
	 ("00000000000000000000000000000000"),	 -- 218	0
	 ("00000000000000000000000000000000"),	 -- 217	0
	 ("00000000000000000000000000000000"),	 -- 216	0
	 ("00000000000000000000000000000000"),	 -- 215	0
	 ("00000000000000000000000000000000"),	 -- 214	0
	 ("00000000000000000000000000000000"),	 -- 213	0
	 ("00000000000000000000000000000000"),	 -- 212	0
	 ("00000000000000000000000000000000"),	 -- 211	0
	 ("00000000000000000000000000000000"),	 -- 210	0
	 ("00000000000000000000000000000000"),	 -- 209	0
	 ("00000000000000000000000000000000"),	 -- 208	0
	 ("00000000000000000000000000000000"),	 -- 207	0
	 ("00000000000000000000000000000000"),	 -- 206	0
	 ("00000000000000000000000000000000"),	 -- 205	0
	 ("00000000000000000000000000000000"),	 -- 204	0
	 ("00000000000000000000000000000000"),	 -- 203	0
	 ("00000000000000000000000000000000"),	 -- 202	0
	 ("00000000000000000000000000000000"),	 -- 201	0
	 ("00000000000000000000000000000000"),	 -- 200	0
	 ("00000000000000000000000000000000"),	 -- 199	0
	 ("00000000000000000000000000000000"),	 -- 198	0
	 ("00000000000000000000000000000000"),	 -- 197	0
	 ("00000000000000000000000000000000"),	 -- 196	0
	 ("00000000000000000000000000000000"),	 -- 195	0
	 ("00000000000000000000000000000000"),	 -- 194	0
	 ("00000000000000000000000000000000"),	 -- 193	0
	 ("00000000000000000000000000000000"),	 -- 192	0
	 ("00000000000000000000000000000000"),	 -- 191	0
	 ("00000000000000000000000000000000"),	 -- 190	0
	 ("00000000000000000000000000000000"),	 -- 189	0
	 ("00000000000000000000000000000000"),	 -- 188	0
	 ("00000000000000000000000000000000"),	 -- 187	0
	 ("00000000000000000000000000000000"),	 -- 186	0
	 ("00000000000000000000000000000000"),	 -- 185	0
	 ("00000000000000000000000000000000"),	 -- 184	0
	 ("00000000000000000000000000000000"),	 -- 183	0
	 ("00000000000000000000000000000000"),	 -- 182	0
	 ("00000000000000000000000000000000"),	 -- 181	0
	 ("00000000000000000000000000000000"),	 -- 180	0
	 ("00000000000000000000000000000000"),	 -- 179	0
	 ("00000000000000000000000000000000"),	 -- 178	0
	 ("00000000000000000000000000000000"),	 -- 177	0
	 ("00000000000000000000000000000000"),	 -- 176	0
	 ("00000000000000000000000000000000"),	 -- 175	0
	 ("00000000000000000000000000000000"),	 -- 174	0
	 ("00000000000000000000000000000000"),	 -- 173	0
	 ("00000000000000000000000000000000"),	 -- 172	0
	 ("00000000000000000000000000000000"),	 -- 171	0
	 ("00000000000000000000000000000000"),	 -- 170	0
	 ("00000000000000000000000000000000"),	 -- 169	0
	 ("00000000000000000000000000000000"),	 -- 168	0
	 ("00000000000000000000000000000000"),	 -- 167	0
	 ("00000000000000000000000000000000"),	 -- 166	0
	 ("00000000000000000000000000000000"),	 -- 165	0
	 ("00000000000000000000000000000000"),	 -- 164	0
	 ("00000000000000000000000000000000"),	 -- 163	0
	 ("00000000000000000000000000000000"),	 -- 162	0
	 ("00000000000000000000000000000000"),	 -- 161	0
	 ("00000000000000000000000000000000"),	 -- 160	0
	 ("00000000000000000000000000000000"),	 -- 159	0
	 ("00000000000000000000000000000000"),	 -- 158	0
	 ("00000000000000000000000000000000"),	 -- 157	0
	 ("00000000000000000000000000000000"),	 -- 156	0
	 ("00000000000000000000000000000000"),	 -- 155	0
	 ("00000000000000000000000000000000"),	 -- 154	0
	 ("00000000000000000000000000000000"),	 -- 153	0
	 ("00000000000000000000000000000000"),	 -- 152	0
	 ("00000000000000000000000000000000"),	 -- 151	0
	 ("00000000000000000000000000000000"),	 -- 150	0
	 ("00000000000000000000000000000000"),	 -- 149	0
	 ("00000000000000000000000000000000"),	 -- 148	0
	 ("00000000000000000000000000000000"),	 -- 147	0
	 ("00000000000000000000000000000000"),	 -- 146	0
	 ("00000000000000000000000000000000"),	 -- 145	0
	 ("00000000000000000000000000000000"),	 -- 144	0
	 ("00000000000000000000000000000000"),	 -- 143	0
	 ("00000000000000000000000000000000"),	 -- 142	0
	 ("00000000000000000000000000000000"),	 -- 141	0
	 ("00000000000000000000000000000000"),	 -- 140	0
	 ("00000000000000000000000000000000"),	 -- 139	0
	 ("00000000000000000000000000000000"),	 -- 138	0
	 ("00000000000000000000000000000000"),	 -- 137	0
	 ("00000000000000000000000000000000"),	 -- 136	0
	 ("00000000000000000000000000000000"),	 -- 135	0
	 ("00000000000000000000000000000000"),	 -- 134	0
	 ("00000000000000000000000000000000"),	 -- 133	0
	 ("00000000000000000000000000000000"),	 -- 132	0
	 ("00000000000000000000000000000000"),	 -- 131	0
	 ("00000000000000000000000000000000"),	 -- 130	0
	 ("00000000000000000000000000000000"),	 -- 129	0
	 ("00000000000000000000000000000000"),	 -- 128	0
	 ("00000000000000000000000000000000"),	 -- 127	0
	 ("00000000000000000000000000000000"),	 -- 126	0
	 ("00000000000000000000000000000000"),	 -- 125	0
	 ("00000000000000000000000000000000"),	 -- 124	0
	 ("00000000000000000000000000000000"),	 -- 123	0
	 ("00000000000000000000000000000000"),	 -- 122	0
	 ("00000000000000000000000000000000"),	 -- 121	0
	 ("00000000000000000000000000000000"),	 -- 120	0
	 ("00000000000000000000000000000000"),	 -- 119	0
	 ("00000000000000000000000000000000"),	 -- 118	0
	 ("00000000000000000000000000000000"),	 -- 117	0
	 ("00000000000000000000000000000000"),	 -- 116	0
	 ("00000000000000000000000000000000"),	 -- 115	0
	 ("00000000000000000000000000000000"),	 -- 114	0
	 ("00000000000000000000000000000000"),	 -- 113	0
	 ("00000000000000000000000000000000"),	 -- 112	0
	 ("00000000000000000000000000000000"),	 -- 111	0
	 ("00000000000000000000000000000000"),	 -- 110	0
	 ("00000000000000000000000000000000"),	 -- 109	0
	 ("00000000000000000000000000000000"),	 -- 108	0
	 ("00000000000000000000000000000000"),	 -- 107	0
	 ("00000000000000000000000000000000"),	 -- 106	0
	 ("00000000000000000000000000000000"),	 -- 105	0
	 ("00000000000000000000000000000000"),	 -- 104	0
	 ("00000000000000000000000000000000"),	 -- 103	0
	 ("00000000000000000000000000000000"),	 -- 102	0
	 ("00000000000000000000000000000000"),	 -- 101	0
	 ("00000000000000000000000000000000"),	 -- 100	0
	 ("00000000000000000000000000000000"),	 -- 99	0
	 ("00000000000000000000000000000000"),	 -- 98	0
	 ("00000000000000000000000000000000"),	 -- 97	0
	 ("00000000000000000000000000000000"),	 -- 96	0
	 ("00000000000000000000000000000000"),	 -- 95	0
	 ("00000000000000000000000000000000"),	 -- 94	0
	 ("00000000000000000000000000000000"),	 -- 93	0
	 ("00000000000000000000000000000000"),	 -- 92	0
	 ("00000000000000000000000000000000"),	 -- 91	0
	 ("00000000000000000000000000000000"),	 -- 90	0
	 ("00000000000000000000000000000000"),	 -- 89	0
	 ("00000000000000000000000000000000"),	 -- 88	0
	 ("00000000000000000000000000000000"),	 -- 87	0
	 ("00000000000000000000000000000000"),	 -- 86	0
	 ("00000000000000000000000000000000"),	 -- 85	0
	 ("00000000000000000000000000000000"),	 -- 84	0
	 ("00000000000000000000000000000000"),	 -- 83	0
	 ("00000000000000000000000000000000"),	 -- 82	0
	 ("00000000000000000000000000000000"),	 -- 81	0
	 ("00000000000000000000000000000000"),	 -- 80	0
	 ("00000000000000000000000000000000"),	 -- 79	0
	 ("00000000000000000000000000000000"),	 -- 78	0
	 ("00000000000000000000000000000000"),	 -- 77	0
	 ("00000000000000000000000000000000"),	 -- 76	0
	 ("00000000000000000000000000000000"),	 -- 75	0
	 ("00000000000000000000000000000000"),	 -- 74	0
	 ("00000000000000000000000000000000"),	 -- 73	0
	 ("00000000000000000000000000000000"),	 -- 72	0
	 ("00000000000000000000000000000000"),	 -- 71	0
	 ("00000000000000000000000000000000"),	 -- 70	0
	 ("00000000000000000000000000000000"),	 -- 69	0
	 ("00000000000000000000000000000000"),	 -- 68	0
	 ("00000000000000000000000000000000"),	 -- 67	0
	 ("00000000000000000000000000000000"),	 -- 66	0
	 ("00000000000000000000000000000000"),	 -- 65	0
	 ("00000000000000000000000000000000"),	 -- 64	0
	 ("00000000000000000000000000000000"),	 -- 63	0
	 ("00000000000000000000000000000000"),	 -- 62	0
	 ("00000000000000000000000000000000"),	 -- 61	0
	 ("00000000000000000000000000000000"),	 -- 60	0
	 ("00000000000000000000000000000000"),	 -- 59	0
	 ("00000000000000000000000000000000"),	 -- 58	0
	 ("00000000000000000000000000000000"),	 -- 57	0
	 ("00000000000000000000000000000000"),	 -- 56	0
	 ("00000000000000000000000000000000"),	 -- 55	0
	 ("00000000000000000000000000000000"),	 -- 54	0
	 ("00000000000000000000000000000000"),	 -- 53	0
	 ("00000000000000000000000000000000"),	 -- 52	0
	 ("00000000000000000000000000000000"),	 -- 51	0
	 ("00000000000000000000000000000000"),	 -- 50	0
	 ("00000000000000000000000000000000"),	 -- 49	0
	 ("00000000000000000000000000000000"),	 -- 48	0
	 ("00000000000000000000000000000000"),	 -- 47	0
	 ("00000000000000000000000000000000"),	 -- 46	0
	 ("00000000000000000000000000000000"),	 -- 45	0
	 ("00000000000000000000000000000000"),	 -- 44	0
	 ("00000000000000000000000000000000"),	 -- 43	0
	 ("00000000000000000000000000000000"),	 -- 42	0
	 ("00000000000000000000000000000000"),	 -- 41	0
	 ("00000000000000000000000000000000"),	 -- 40	0
	 ("00000000000000000000000000000000"),	 -- 39	0
	 ("00000000000000000000000000000000"),	 -- 38	0
	 ("00000000000000000000000000000000"),	 -- 37	0
	 ("00000000000000000000000000000000"),	 -- 36	0
	 ("00000000000000000000000000000000"),	 -- 35	0
	 ("00000000000000000000000000000000"),	 -- 34	0
	 ("00000000000000000000000000000000"),	 -- 33	0
	 ("00000000000000000000000000000000"),	 -- 32	0
	 ("00000000000000000000000000000000"),	 -- 31	0
	 ("00000000000000000000000000000000"),	 -- 30	0
	 ("00000000000000000000000000000000"),	 -- 29	0
	 ("00000000000000000000000000000000"),	 -- 28	0
	 ("00000000000000000000000000000000"),	 -- 27	0
	 ("00000000000000000000000000000000"),	 -- 26	0
	 ("00000000000000000000000000000000"),	 -- 25	0
	 ("00000000000000000000000000000000"),	 -- 24	0
	 ("00000000000000000000000000000000"),	 -- 23	0
	 ("00000000000000000000000000000000"),	 -- 22	0
	 ("00000000000000000000000000000000"),	 -- 21	0
	 ("00000000000000000000000000000000"),	 -- 20	0
	 ("00000000000000000000000000000000"),	 -- 19	0
	 ("00000000000000000000000000000000"),	 -- 18	0
	 ("00000000000000000000000000000000"),	 -- 17	0
	 ("00000000000000000000000000000000"),	 -- 16	0
	 ("00000000000000000000000000000000"),	 -- 15	0
	 ("00000000000000000000000000000000"),	 -- 14	0
	 ("00000000000000000000000000000000"),	 -- 13	0
	 ("00000000000000000000000000000000"),	 -- 12	0
	 ("00000000000000000000000000000000"),	 -- 11	0
	 ("00000000000000000000000000000000"),	 -- 10	0
	 ("00000000000000000000000000000000"),	 -- 9	0
	 ("00000000000000000000000000000000"),	 -- 8	0
	 ("00000000000000000000000000000000"),	 -- 7	0
	 ("00000000000000000000000000000000"),	 -- 6	0
	 ("00000000000000000000000000000000"),	 -- 5	0
	 ("00000000000000000000000000000000"),	 -- 4	0
	 ("00000000000000000000000000000000"),	 -- 3	0
	 ("00000000000000000000000000000011"),	 -- 2	3
	 ("00000000000000000000000000000100"),	 -- 1	4
	 ("00000000000000000000000000000110"));	 -- 0	6


begin 
       process (clk) 
       begin 
              if (clk'event and clk = '1') then 
                  if (we_0 = '1') then 
                        RAM(conv_integer(address_0)) <= data_in_0; 
                        data_out_0 <= RAM(conv_integer(read_a)); 
                  elsif (oe_0 = '1') then 
                        data_out_0 <= RAM(conv_integer(read_a)); 
                  end if; 
                  read_a <= address_0; 
             end if; 
       end process; 
       process (clk) 
       begin 
              if (clk'event and clk = '1') then 
                  if (we_1 = '1') then 
                        RAM(conv_integer(address_1)) <= data_in_1; 
                        data_out_1 <= RAM(conv_integer(read_b)); 
                  elsif (oe_1 = '1') then 
                        data_out_1 <= RAM(conv_integer(read_b)); 
                  end if; 
                  read_b <= address_1; 
             end if; 
       end process; 
end rtl; 

