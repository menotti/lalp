library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 
entity vecsum is 
	port (
		\init\	: in	std_logic;
		\done\	: out	std_logic;
		\out_19\	: out	std_logic_vector(31 downto 0);
		\clk\	: in	std_logic;
		\reset\	: in	std_logic;
		\clear\	: in	std_logic
	);
end vecsum; 

architecture behavior of vecsum is 

component add_op_s 
generic ( 
        w_in1	: integer := 8; 
        w_in2	: integer := 8; 
        w_out	: integer := 16 
); 
port ( 
        I0          : in	std_logic_vector(w_in1-1 downto 0); 
        I1          : in	std_logic_vector(w_in2-1 downto 0); 
        O0          : out	std_logic_vector(w_out-1 downto 0) 
); 
end component; 

component block_ram 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_x 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component block_ram_y 
generic ( 
        data_width          : integer := 8; 
        address_width	: integer := 8 
); 
port ( 
        clk                 : in	std_logic; 
        we                  : in	std_logic := '0'; 
        oe                  : in	std_logic := '1'; 
        address             : in	std_logic_vector(address_width-1 downto 0); 
        data_in             : in	std_logic_vector(data_width-1 downto 0) := (others => '0'); 
        data_out            : out	std_logic_vector(data_width-1 downto 0) 
); 
end component; 

component counter 
generic (
        bits		: integer := 8;
        steps		: integer := 1;
        increment           : integer := 1;
        down                : integer := 0;
        condition           : integer := 0
);
port (
        input		: in	std_logic_vector(bits-1 downto 0);
        termination         : in	std_logic_vector(bits-1 downto 0);
        clk                 : in	std_logic;
        clk_en		: in	std_logic := '1';
        reset		: in	std_logic;
        load		: in	std_logic := '0';
        step		: out	std_logic;
        done		: out	std_logic;
        output		: out	std_logic_vector(bits-1 downto 0)
); 
end component; 

component delay_op 
generic ( 
        bits        : integer := 8; 
        delay       : integer := 1 
); 
port ( 
        a		: in	std_logic_vector(bits-1 downto 0); 
        clk		: in	std_logic; 
        reset	: in	std_logic; 
        a_delayed	: out	std_logic_vector(bits-1 downto 0) := (others=>'0') 
); 
end component; 

signal s2	: std_logic_vector(31 downto 0); 
signal s3	: std_logic_vector(31 downto 0); 
signal s4	: std_logic_vector(31 downto 0); 
signal s5	: std_logic_vector(31 downto 0); 
signal s6	: std_logic_vector(31 downto 0); 
signal s7	: std_logic_vector(31 downto 0); 
signal s8	: std_logic_vector(31 downto 0); 
signal s9	: std_logic; 
signal s10	: std_logic_vector(0 downto 0); 
signal s11	: std_logic; 
signal s12	: std_logic; 
signal s13	: std_logic_vector(0 downto 0); 
signal s14	: std_logic_vector(31 downto 0); 

begin 

\i\: counter
generic map ( 
	bits => 32,
	condition => 0,
	down => 0,
	increment => 1,
	steps => 1
)
port map ( 
	clk => \clk\,
	clk_en => s11,
	done => s12,
	input => s7,
	output => s2,
	reset => \reset\,
	step => s9,
	termination => s6
);

\z\: block_ram
generic map ( 
	address_width => 11,
	data_width => 32
)
port map ( 
	address(10 downto 0) => s8(10 downto 0),
	clk => \clk\,
	data_in => s3,
	data_out => s14,
	we => s10(0)
);

\x_add_op_s_y\: add_op_s
generic map ( 
	w_in1 => 32,
	w_in2 => 32,
	w_out => 32
)
port map ( 
	I0 => s4,
	I1 => s5,
	O0 => s3
);

\x\: block_ram_x
generic map ( 
	address_width => 11,
	data_width => 32
)
port map ( 
	address(10 downto 0) => s2(10 downto 0),
	clk => \clk\,
	data_out => s4
);

\y\: block_ram_y
generic map ( 
	address_width => 11,
	data_width => 32
)
port map ( 
	address(10 downto 0) => s2(10 downto 0),
	clk => \clk\,
	data_out => s5
);

\dly_16\: delay_op
generic map ( 
	bits => 32,
	delay => 2
)
port map ( 
	a => s2,
	a_delayed => s8,
	clk => \clk\,
	reset => \reset\
);

\dly_17\: delay_op
generic map ( 
	bits => 1,
	delay => 2
)
port map ( 
	a(0) => s9,
	a_delayed => s10,
	clk => \clk\,
	reset => \reset\
);

\dly_18\: delay_op
generic map ( 
	bits => 1,
	delay => 4
)
port map ( 
	a(0) => s12,
	a_delayed => s13,
	clk => \clk\,
	reset => \reset\
);

s11 <= \init\;
\done\ <= s13(0);
s6 <= conv_std_logic_vector(2048, 32);
s7 <= conv_std_logic_vector(0, 32);
\out_19\ <= s14;
end behavior; 