library IEEE; 
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 
entity accumulation is 
	port (
		\init\	: in	std_logic;
		\done\	: out	std_logic;
		\clk\	: in	std_logic;
		\reset\	: in	std_logic;
		\clear\	: in	std_logic
	);
end accumulation; 

architecture behavior of accumulation is 


begin 

end behavior; 