--
-- Copyright (c) 2010 Ricardo Menotti, All Rights Reserved.
--
-- Permission to use, copy, modify, and distribute this software and its
-- documentation for NON-COMERCIAL purposes and without fee is hereby granted 
-- provided that this copyright notice appears in all copies.
--
-- RICARDO MENOTTI MAKES NO REPRESENTATIONS OR WARRANTIES ABOUT THE SUITABILITY
-- OF THE SOFTWARE, EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE, OR
-- NON-INFRINGEMENT. RICARDO MENOTTI SHALL NOT BE LIABLE FOR ANY DAMAGES
-- SUFFERED BY LICENSEE AS A RESULT OF USING, MODIFYING OR DISTRIBUTING THIS
-- SOFTWARE OR ITS DERIVATIVES.
--
-- Generated at Tue May 10 19:39:40 BRT 2011
--

-- IEEE Libraries --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity block_ram_v is
generic(
	data_width : integer := 8;
	address_width : integer := 8
);
port(
	data_in : in std_logic_vector(data_width-1 downto 0) := (others => '0');
	address : in std_logic_vector(address_width-1 downto 0);
	we: in std_logic := '0';
	oe: in std_logic := '1';
	clk : in std_logic;
	data_out : out std_logic_vector(data_width-1 downto 0));
end block_ram_v;

architecture rtl of block_ram_v is

constant mem_depth : integer := 2**address_width;
type ram_type is array (mem_depth-1 downto 0)
of std_logic_vector (data_width-1 downto 0);

signal read_a : std_logic_vector(address_width-1 downto 0);
signal RAM : ram_type := ram_type'(
	 ("00000000000000000000001100100000"),	 -- 2047	800
	 ("00000000000000000000000000000111"),	 -- 2046	7
	 ("00000000000000000000000000000110"),	 -- 2045	6
	 ("00000000000000000000000000000101"),	 -- 2044	5
	 ("00000000000000000000000000000100"),	 -- 2043	4
	 ("00000000000000000000000000000011"),	 -- 2042	3
	 ("00000000000000000000000000000010"),	 -- 2041	2
	 ("00000000000000000000000000000001"),	 -- 2040	1
	 ("00000000000000000000000000001000"),	 -- 2039	8
	 ("00000000000000000000000000000111"),	 -- 2038	7
	 ("00000000000000000000000000000110"),	 -- 2037	6
	 ("00000000000000000000000000000101"),	 -- 2036	5
	 ("00000000000000000000000000000100"),	 -- 2035	4
	 ("00000000000000000000000000000011"),	 -- 2034	3
	 ("00000000000000000000000000000010"),	 -- 2033	2
	 ("00000000000000000000000000000001"),	 -- 2032	1
	 ("00000000000000000000000000001000"),	 -- 2031	8
	 ("00000000000000000000000000000111"),	 -- 2030	7
	 ("00000000000000000000000000000110"),	 -- 2029	6
	 ("00000000000000000000000000000101"),	 -- 2028	5
	 ("00000000000000000000000000000100"),	 -- 2027	4
	 ("00000000000000000000000000000011"),	 -- 2026	3
	 ("00000000000000000000000000000010"),	 -- 2025	2
	 ("00000000000000000000000000000001"),	 -- 2024	1
	 ("00000000000000000000000000001000"),	 -- 2023	8
	 ("00000000000000000000000000000111"),	 -- 2022	7
	 ("00000000000000000000000000000110"),	 -- 2021	6
	 ("00000000000000000000000000000101"),	 -- 2020	5
	 ("00000000000000000000000000000100"),	 -- 2019	4
	 ("00000000000000000000000000000011"),	 -- 2018	3
	 ("00000000000000000000000000000010"),	 -- 2017	2
	 ("00000000000000000000000000000001"),	 -- 2016	1
	 ("00000000000000000000000000001000"),	 -- 2015	8
	 ("00000000000000000000000000000111"),	 -- 2014	7
	 ("00000000000000000000000000000110"),	 -- 2013	6
	 ("00000000000000000000000000000101"),	 -- 2012	5
	 ("00000000000000000000000000000100"),	 -- 2011	4
	 ("00000000000000000000000000000011"),	 -- 2010	3
	 ("00000000000000000000000000000010"),	 -- 2009	2
	 ("00000000000000000000000000000001"),	 -- 2008	1
	 ("00000000000000000000000000001000"),	 -- 2007	8
	 ("00000000000000000000000000000111"),	 -- 2006	7
	 ("00000000000000000000000000000110"),	 -- 2005	6
	 ("00000000000000000000000000000101"),	 -- 2004	5
	 ("00000000000000000000000000000100"),	 -- 2003	4
	 ("00000000000000000000000000000011"),	 -- 2002	3
	 ("00000000000000000000000000000010"),	 -- 2001	2
	 ("00000000000000000000000000000001"),	 -- 2000	1
	 ("00000000000000000000000000001000"),	 -- 1999	8
	 ("00000000000000000000000000000111"),	 -- 1998	7
	 ("00000000000000000000000000000110"),	 -- 1997	6
	 ("00000000000000000000000000000101"),	 -- 1996	5
	 ("00000000000000000000000000000100"),	 -- 1995	4
	 ("00000000000000000000000000000011"),	 -- 1994	3
	 ("00000000000000000000000000000010"),	 -- 1993	2
	 ("00000000000000000000000000000001"),	 -- 1992	1
	 ("00000000000000000000000000001000"),	 -- 1991	8
	 ("00000000000000000000000000000111"),	 -- 1990	7
	 ("00000000000000000000000000000110"),	 -- 1989	6
	 ("00000000000000000000000000000101"),	 -- 1988	5
	 ("00000000000000000000000000000100"),	 -- 1987	4
	 ("00000000000000000000000000000011"),	 -- 1986	3
	 ("00000000000000000000000000000010"),	 -- 1985	2
	 ("00000000000000000000000000000001"),	 -- 1984	1
	 ("00000000000000000000000000001000"),	 -- 1983	8
	 ("00000000000000000000000000000111"),	 -- 1982	7
	 ("00000000000000000000000000000110"),	 -- 1981	6
	 ("00000000000000000000000000000101"),	 -- 1980	5
	 ("00000000000000000000000000000100"),	 -- 1979	4
	 ("00000000000000000000000000000011"),	 -- 1978	3
	 ("00000000000000000000000000000010"),	 -- 1977	2
	 ("00000000000000000000000000000001"),	 -- 1976	1
	 ("00000000000000000000000000001000"),	 -- 1975	8
	 ("00000000000000000000000000000111"),	 -- 1974	7
	 ("00000000000000000000000000000110"),	 -- 1973	6
	 ("00000000000000000000000000000101"),	 -- 1972	5
	 ("00000000000000000000000000000100"),	 -- 1971	4
	 ("00000000000000000000000000000011"),	 -- 1970	3
	 ("00000000000000000000000000000010"),	 -- 1969	2
	 ("00000000000000000000000000000001"),	 -- 1968	1
	 ("00000000000000000000000000001000"),	 -- 1967	8
	 ("00000000000000000000000000000111"),	 -- 1966	7
	 ("00000000000000000000000000000110"),	 -- 1965	6
	 ("00000000000000000000000000000101"),	 -- 1964	5
	 ("00000000000000000000000000000100"),	 -- 1963	4
	 ("00000000000000000000000000000011"),	 -- 1962	3
	 ("00000000000000000000000000000010"),	 -- 1961	2
	 ("00000000000000000000000000000001"),	 -- 1960	1
	 ("00000000000000000000000000001000"),	 -- 1959	8
	 ("00000000000000000000000000000111"),	 -- 1958	7
	 ("00000000000000000000000000000110"),	 -- 1957	6
	 ("00000000000000000000000000000101"),	 -- 1956	5
	 ("00000000000000000000000000000100"),	 -- 1955	4
	 ("00000000000000000000000000000011"),	 -- 1954	3
	 ("00000000000000000000000000000010"),	 -- 1953	2
	 ("00000000000000000000000000000001"),	 -- 1952	1
	 ("00000000000000000000000000001000"),	 -- 1951	8
	 ("00000000000000000000000000000111"),	 -- 1950	7
	 ("00000000000000000000000000000110"),	 -- 1949	6
	 ("00000000000000000000000000000101"),	 -- 1948	5
	 ("00000000000000000000000000000100"),	 -- 1947	4
	 ("00000000000000000000000000000011"),	 -- 1946	3
	 ("00000000000000000000000000000010"),	 -- 1945	2
	 ("00000000000000000000000000000001"),	 -- 1944	1
	 ("00000000000000000000000000001000"),	 -- 1943	8
	 ("00000000000000000000000000000111"),	 -- 1942	7
	 ("00000000000000000000000000000110"),	 -- 1941	6
	 ("00000000000000000000000000000101"),	 -- 1940	5
	 ("00000000000000000000000000000100"),	 -- 1939	4
	 ("00000000000000000000000000000011"),	 -- 1938	3
	 ("00000000000000000000000000000010"),	 -- 1937	2
	 ("00000000000000000000000000000001"),	 -- 1936	1
	 ("00000000000000000000000000001000"),	 -- 1935	8
	 ("00000000000000000000000000000111"),	 -- 1934	7
	 ("00000000000000000000000000000110"),	 -- 1933	6
	 ("00000000000000000000000000000101"),	 -- 1932	5
	 ("00000000000000000000000000000100"),	 -- 1931	4
	 ("00000000000000000000000000000011"),	 -- 1930	3
	 ("00000000000000000000000000000010"),	 -- 1929	2
	 ("00000000000000000000000000000001"),	 -- 1928	1
	 ("00000000000000000000000000001000"),	 -- 1927	8
	 ("00000000000000000000000000000111"),	 -- 1926	7
	 ("00000000000000000000000000000110"),	 -- 1925	6
	 ("00000000000000000000000000000101"),	 -- 1924	5
	 ("00000000000000000000000000000100"),	 -- 1923	4
	 ("00000000000000000000000000000011"),	 -- 1922	3
	 ("00000000000000000000000000000010"),	 -- 1921	2
	 ("00000000000000000000000000000001"),	 -- 1920	1
	 ("00000000000000000000000000001000"),	 -- 1919	8
	 ("00000000000000000000000000000111"),	 -- 1918	7
	 ("00000000000000000000000000000110"),	 -- 1917	6
	 ("00000000000000000000000000000101"),	 -- 1916	5
	 ("00000000000000000000000000000100"),	 -- 1915	4
	 ("00000000000000000000000000000011"),	 -- 1914	3
	 ("00000000000000000000000000000010"),	 -- 1913	2
	 ("00000000000000000000000000000001"),	 -- 1912	1
	 ("00000000000000000000000000001000"),	 -- 1911	8
	 ("00000000000000000000000000000111"),	 -- 1910	7
	 ("00000000000000000000000000000110"),	 -- 1909	6
	 ("00000000000000000000000000000101"),	 -- 1908	5
	 ("00000000000000000000000000000100"),	 -- 1907	4
	 ("00000000000000000000000000000011"),	 -- 1906	3
	 ("00000000000000000000000000000010"),	 -- 1905	2
	 ("00000000000000000000000000000001"),	 -- 1904	1
	 ("00000000000000000000000000001000"),	 -- 1903	8
	 ("00000000000000000000000000000111"),	 -- 1902	7
	 ("00000000000000000000000000000110"),	 -- 1901	6
	 ("00000000000000000000000000000101"),	 -- 1900	5
	 ("00000000000000000000000000000100"),	 -- 1899	4
	 ("00000000000000000000000000000011"),	 -- 1898	3
	 ("00000000000000000000000000000010"),	 -- 1897	2
	 ("00000000000000000000000000000001"),	 -- 1896	1
	 ("00000000000000000000000000001000"),	 -- 1895	8
	 ("00000000000000000000000000000111"),	 -- 1894	7
	 ("00000000000000000000000000000110"),	 -- 1893	6
	 ("00000000000000000000000000000101"),	 -- 1892	5
	 ("00000000000000000000000000000100"),	 -- 1891	4
	 ("00000000000000000000000000000011"),	 -- 1890	3
	 ("00000000000000000000000000000010"),	 -- 1889	2
	 ("00000000000000000000000000000001"),	 -- 1888	1
	 ("00000000000000000000000000001000"),	 -- 1887	8
	 ("00000000000000000000000000000111"),	 -- 1886	7
	 ("00000000000000000000000000000110"),	 -- 1885	6
	 ("00000000000000000000000000000101"),	 -- 1884	5
	 ("00000000000000000000000000000100"),	 -- 1883	4
	 ("00000000000000000000000000000011"),	 -- 1882	3
	 ("00000000000000000000000000000010"),	 -- 1881	2
	 ("00000000000000000000000000000001"),	 -- 1880	1
	 ("00000000000000000000000000001000"),	 -- 1879	8
	 ("00000000000000000000000000000111"),	 -- 1878	7
	 ("00000000000000000000000000000110"),	 -- 1877	6
	 ("00000000000000000000000000000101"),	 -- 1876	5
	 ("00000000000000000000000000000100"),	 -- 1875	4
	 ("00000000000000000000000000000011"),	 -- 1874	3
	 ("00000000000000000000000000000010"),	 -- 1873	2
	 ("00000000000000000000000000000001"),	 -- 1872	1
	 ("00000000000000000000000000001000"),	 -- 1871	8
	 ("00000000000000000000000000000111"),	 -- 1870	7
	 ("00000000000000000000000000000110"),	 -- 1869	6
	 ("00000000000000000000000000000101"),	 -- 1868	5
	 ("00000000000000000000000000000100"),	 -- 1867	4
	 ("00000000000000000000000000000011"),	 -- 1866	3
	 ("00000000000000000000000000000010"),	 -- 1865	2
	 ("00000000000000000000000000000001"),	 -- 1864	1
	 ("00000000000000000000000000001000"),	 -- 1863	8
	 ("00000000000000000000000000000111"),	 -- 1862	7
	 ("00000000000000000000000000000110"),	 -- 1861	6
	 ("00000000000000000000000000000101"),	 -- 1860	5
	 ("00000000000000000000000000000100"),	 -- 1859	4
	 ("00000000000000000000000000000011"),	 -- 1858	3
	 ("00000000000000000000000000000010"),	 -- 1857	2
	 ("00000000000000000000000000000001"),	 -- 1856	1
	 ("00000000000000000000000000001000"),	 -- 1855	8
	 ("00000000000000000000000000000111"),	 -- 1854	7
	 ("00000000000000000000000000000110"),	 -- 1853	6
	 ("00000000000000000000000000000101"),	 -- 1852	5
	 ("00000000000000000000000000000100"),	 -- 1851	4
	 ("00000000000000000000000000000011"),	 -- 1850	3
	 ("00000000000000000000000000000010"),	 -- 1849	2
	 ("00000000000000000000000000000001"),	 -- 1848	1
	 ("00000000000000000000000000001000"),	 -- 1847	8
	 ("00000000000000000000000000000111"),	 -- 1846	7
	 ("00000000000000000000000000000110"),	 -- 1845	6
	 ("00000000000000000000000000000101"),	 -- 1844	5
	 ("00000000000000000000000000000100"),	 -- 1843	4
	 ("00000000000000000000000000000011"),	 -- 1842	3
	 ("00000000000000000000000000000010"),	 -- 1841	2
	 ("00000000000000000000000000000001"),	 -- 1840	1
	 ("00000000000000000000000000001000"),	 -- 1839	8
	 ("00000000000000000000000000000111"),	 -- 1838	7
	 ("00000000000000000000000000000110"),	 -- 1837	6
	 ("00000000000000000000000000000101"),	 -- 1836	5
	 ("00000000000000000000000000000100"),	 -- 1835	4
	 ("00000000000000000000000000000011"),	 -- 1834	3
	 ("00000000000000000000000000000010"),	 -- 1833	2
	 ("00000000000000000000000000000001"),	 -- 1832	1
	 ("00000000000000000000000000001000"),	 -- 1831	8
	 ("00000000000000000000000000000111"),	 -- 1830	7
	 ("00000000000000000000000000000110"),	 -- 1829	6
	 ("00000000000000000000000000000101"),	 -- 1828	5
	 ("00000000000000000000000000000100"),	 -- 1827	4
	 ("00000000000000000000000000000011"),	 -- 1826	3
	 ("00000000000000000000000000000010"),	 -- 1825	2
	 ("00000000000000000000000000000001"),	 -- 1824	1
	 ("00000000000000000000000000001000"),	 -- 1823	8
	 ("00000000000000000000000000000111"),	 -- 1822	7
	 ("00000000000000000000000000000110"),	 -- 1821	6
	 ("00000000000000000000000000000101"),	 -- 1820	5
	 ("00000000000000000000000000000100"),	 -- 1819	4
	 ("00000000000000000000000000000011"),	 -- 1818	3
	 ("00000000000000000000000000000010"),	 -- 1817	2
	 ("00000000000000000000000000000001"),	 -- 1816	1
	 ("00000000000000000000000000001000"),	 -- 1815	8
	 ("00000000000000000000000000000111"),	 -- 1814	7
	 ("00000000000000000000000000000110"),	 -- 1813	6
	 ("00000000000000000000000000000101"),	 -- 1812	5
	 ("00000000000000000000000000000100"),	 -- 1811	4
	 ("00000000000000000000000000000011"),	 -- 1810	3
	 ("00000000000000000000000000000010"),	 -- 1809	2
	 ("00000000000000000000000000000001"),	 -- 1808	1
	 ("00000000000000000000000000001000"),	 -- 1807	8
	 ("00000000000000000000000000000111"),	 -- 1806	7
	 ("00000000000000000000000000000110"),	 -- 1805	6
	 ("00000000000000000000000000000101"),	 -- 1804	5
	 ("00000000000000000000000000000100"),	 -- 1803	4
	 ("00000000000000000000000000000011"),	 -- 1802	3
	 ("00000000000000000000000000000010"),	 -- 1801	2
	 ("00000000000000000000000000000001"),	 -- 1800	1
	 ("00000000000000000000000000001000"),	 -- 1799	8
	 ("00000000000000000000000000000111"),	 -- 1798	7
	 ("00000000000000000000000000000110"),	 -- 1797	6
	 ("00000000000000000000000000000101"),	 -- 1796	5
	 ("00000000000000000000000000000100"),	 -- 1795	4
	 ("00000000000000000000000000000011"),	 -- 1794	3
	 ("00000000000000000000000000000010"),	 -- 1793	2
	 ("00000000000000000000000000000001"),	 -- 1792	1
	 ("00000000000000000000000000001000"),	 -- 1791	8
	 ("00000000000000000000000000000111"),	 -- 1790	7
	 ("00000000000000000000000000000110"),	 -- 1789	6
	 ("00000000000000000000000000000101"),	 -- 1788	5
	 ("00000000000000000000000000000100"),	 -- 1787	4
	 ("00000000000000000000000000000011"),	 -- 1786	3
	 ("00000000000000000000000000000010"),	 -- 1785	2
	 ("00000000000000000000000000000001"),	 -- 1784	1
	 ("00000000000000000000000000001000"),	 -- 1783	8
	 ("00000000000000000000000000000111"),	 -- 1782	7
	 ("00000000000000000000000000000110"),	 -- 1781	6
	 ("00000000000000000000000000000101"),	 -- 1780	5
	 ("00000000000000000000000000000100"),	 -- 1779	4
	 ("00000000000000000000000000000011"),	 -- 1778	3
	 ("00000000000000000000000000000010"),	 -- 1777	2
	 ("00000000000000000000000000000001"),	 -- 1776	1
	 ("00000000000000000000000000001000"),	 -- 1775	8
	 ("00000000000000000000000000000111"),	 -- 1774	7
	 ("00000000000000000000000000000110"),	 -- 1773	6
	 ("00000000000000000000000000000101"),	 -- 1772	5
	 ("00000000000000000000000000000100"),	 -- 1771	4
	 ("00000000000000000000000000000011"),	 -- 1770	3
	 ("00000000000000000000000000000010"),	 -- 1769	2
	 ("00000000000000000000000000000001"),	 -- 1768	1
	 ("00000000000000000000000000001000"),	 -- 1767	8
	 ("00000000000000000000000000000111"),	 -- 1766	7
	 ("00000000000000000000000000000110"),	 -- 1765	6
	 ("00000000000000000000000000000101"),	 -- 1764	5
	 ("00000000000000000000000000000100"),	 -- 1763	4
	 ("00000000000000000000000000000011"),	 -- 1762	3
	 ("00000000000000000000000000000010"),	 -- 1761	2
	 ("00000000000000000000000000000001"),	 -- 1760	1
	 ("00000000000000000000000000001000"),	 -- 1759	8
	 ("00000000000000000000000000000111"),	 -- 1758	7
	 ("00000000000000000000000000000110"),	 -- 1757	6
	 ("00000000000000000000000000000101"),	 -- 1756	5
	 ("00000000000000000000000000000100"),	 -- 1755	4
	 ("00000000000000000000000000000011"),	 -- 1754	3
	 ("00000000000000000000000000000010"),	 -- 1753	2
	 ("00000000000000000000000000000001"),	 -- 1752	1
	 ("00000000000000000000000000001000"),	 -- 1751	8
	 ("00000000000000000000000000000111"),	 -- 1750	7
	 ("00000000000000000000000000000110"),	 -- 1749	6
	 ("00000000000000000000000000000101"),	 -- 1748	5
	 ("00000000000000000000000000000100"),	 -- 1747	4
	 ("00000000000000000000000000000011"),	 -- 1746	3
	 ("00000000000000000000000000000010"),	 -- 1745	2
	 ("00000000000000000000000000000001"),	 -- 1744	1
	 ("00000000000000000000000000001000"),	 -- 1743	8
	 ("00000000000000000000000000000111"),	 -- 1742	7
	 ("00000000000000000000000000000110"),	 -- 1741	6
	 ("00000000000000000000000000000101"),	 -- 1740	5
	 ("00000000000000000000000000000100"),	 -- 1739	4
	 ("00000000000000000000000000000011"),	 -- 1738	3
	 ("00000000000000000000000000000010"),	 -- 1737	2
	 ("00000000000000000000000000000001"),	 -- 1736	1
	 ("00000000000000000000000000001000"),	 -- 1735	8
	 ("00000000000000000000000000000111"),	 -- 1734	7
	 ("00000000000000000000000000000110"),	 -- 1733	6
	 ("00000000000000000000000000000101"),	 -- 1732	5
	 ("00000000000000000000000000000100"),	 -- 1731	4
	 ("00000000000000000000000000000011"),	 -- 1730	3
	 ("00000000000000000000000000000010"),	 -- 1729	2
	 ("00000000000000000000000000000001"),	 -- 1728	1
	 ("00000000000000000000000000001000"),	 -- 1727	8
	 ("00000000000000000000000000000111"),	 -- 1726	7
	 ("00000000000000000000000000000110"),	 -- 1725	6
	 ("00000000000000000000000000000101"),	 -- 1724	5
	 ("00000000000000000000000000000100"),	 -- 1723	4
	 ("00000000000000000000000000000011"),	 -- 1722	3
	 ("00000000000000000000000000000010"),	 -- 1721	2
	 ("00000000000000000000000000000001"),	 -- 1720	1
	 ("00000000000000000000000000001000"),	 -- 1719	8
	 ("00000000000000000000000000000111"),	 -- 1718	7
	 ("00000000000000000000000000000110"),	 -- 1717	6
	 ("00000000000000000000000000000101"),	 -- 1716	5
	 ("00000000000000000000000000000100"),	 -- 1715	4
	 ("00000000000000000000000000000011"),	 -- 1714	3
	 ("00000000000000000000000000000010"),	 -- 1713	2
	 ("00000000000000000000000000000001"),	 -- 1712	1
	 ("00000000000000000000000000001000"),	 -- 1711	8
	 ("00000000000000000000000000000111"),	 -- 1710	7
	 ("00000000000000000000000000000110"),	 -- 1709	6
	 ("00000000000000000000000000000101"),	 -- 1708	5
	 ("00000000000000000000000000000100"),	 -- 1707	4
	 ("00000000000000000000000000000011"),	 -- 1706	3
	 ("00000000000000000000000000000010"),	 -- 1705	2
	 ("00000000000000000000000000000001"),	 -- 1704	1
	 ("00000000000000000000000000001000"),	 -- 1703	8
	 ("00000000000000000000000000000111"),	 -- 1702	7
	 ("00000000000000000000000000000110"),	 -- 1701	6
	 ("00000000000000000000000000000101"),	 -- 1700	5
	 ("00000000000000000000000000000100"),	 -- 1699	4
	 ("00000000000000000000000000000011"),	 -- 1698	3
	 ("00000000000000000000000000000010"),	 -- 1697	2
	 ("00000000000000000000000000000001"),	 -- 1696	1
	 ("00000000000000000000000000001000"),	 -- 1695	8
	 ("00000000000000000000000000000111"),	 -- 1694	7
	 ("00000000000000000000000000000110"),	 -- 1693	6
	 ("00000000000000000000000000000101"),	 -- 1692	5
	 ("00000000000000000000000000000100"),	 -- 1691	4
	 ("00000000000000000000000000000011"),	 -- 1690	3
	 ("00000000000000000000000000000010"),	 -- 1689	2
	 ("00000000000000000000000000000001"),	 -- 1688	1
	 ("00000000000000000000000000001000"),	 -- 1687	8
	 ("00000000000000000000000000000111"),	 -- 1686	7
	 ("00000000000000000000000000000110"),	 -- 1685	6
	 ("00000000000000000000000000000101"),	 -- 1684	5
	 ("00000000000000000000000000000100"),	 -- 1683	4
	 ("00000000000000000000000000000011"),	 -- 1682	3
	 ("00000000000000000000000000000010"),	 -- 1681	2
	 ("00000000000000000000000000000001"),	 -- 1680	1
	 ("00000000000000000000000000001000"),	 -- 1679	8
	 ("00000000000000000000000000000111"),	 -- 1678	7
	 ("00000000000000000000000000000110"),	 -- 1677	6
	 ("00000000000000000000000000000101"),	 -- 1676	5
	 ("00000000000000000000000000000100"),	 -- 1675	4
	 ("00000000000000000000000000000011"),	 -- 1674	3
	 ("00000000000000000000000000000010"),	 -- 1673	2
	 ("00000000000000000000000000000001"),	 -- 1672	1
	 ("00000000000000000000000000001000"),	 -- 1671	8
	 ("00000000000000000000000000000111"),	 -- 1670	7
	 ("00000000000000000000000000000110"),	 -- 1669	6
	 ("00000000000000000000000000000101"),	 -- 1668	5
	 ("00000000000000000000000000000100"),	 -- 1667	4
	 ("00000000000000000000000000000011"),	 -- 1666	3
	 ("00000000000000000000000000000010"),	 -- 1665	2
	 ("00000000000000000000000000000001"),	 -- 1664	1
	 ("00000000000000000000000000001000"),	 -- 1663	8
	 ("00000000000000000000000000000111"),	 -- 1662	7
	 ("00000000000000000000000000000110"),	 -- 1661	6
	 ("00000000000000000000000000000101"),	 -- 1660	5
	 ("00000000000000000000000000000100"),	 -- 1659	4
	 ("00000000000000000000000000000011"),	 -- 1658	3
	 ("00000000000000000000000000000010"),	 -- 1657	2
	 ("00000000000000000000000000000001"),	 -- 1656	1
	 ("00000000000000000000000000001000"),	 -- 1655	8
	 ("00000000000000000000000000000111"),	 -- 1654	7
	 ("00000000000000000000000000000110"),	 -- 1653	6
	 ("00000000000000000000000000000101"),	 -- 1652	5
	 ("00000000000000000000000000000100"),	 -- 1651	4
	 ("00000000000000000000000000000011"),	 -- 1650	3
	 ("00000000000000000000000000000010"),	 -- 1649	2
	 ("00000000000000000000000000000001"),	 -- 1648	1
	 ("00000000000000000000000000001000"),	 -- 1647	8
	 ("00000000000000000000000000000111"),	 -- 1646	7
	 ("00000000000000000000000000000110"),	 -- 1645	6
	 ("00000000000000000000000000000101"),	 -- 1644	5
	 ("00000000000000000000000000000100"),	 -- 1643	4
	 ("00000000000000000000000000000011"),	 -- 1642	3
	 ("00000000000000000000000000000010"),	 -- 1641	2
	 ("00000000000000000000000000000001"),	 -- 1640	1
	 ("00000000000000000000000000001000"),	 -- 1639	8
	 ("00000000000000000000000000000111"),	 -- 1638	7
	 ("00000000000000000000000000000110"),	 -- 1637	6
	 ("00000000000000000000000000000101"),	 -- 1636	5
	 ("00000000000000000000000000000100"),	 -- 1635	4
	 ("00000000000000000000000000000011"),	 -- 1634	3
	 ("00000000000000000000000000000010"),	 -- 1633	2
	 ("00000000000000000000000000000001"),	 -- 1632	1
	 ("00000000000000000000000000001000"),	 -- 1631	8
	 ("00000000000000000000000000000111"),	 -- 1630	7
	 ("00000000000000000000000000000110"),	 -- 1629	6
	 ("00000000000000000000000000000101"),	 -- 1628	5
	 ("00000000000000000000000000000100"),	 -- 1627	4
	 ("00000000000000000000000000000011"),	 -- 1626	3
	 ("00000000000000000000000000000010"),	 -- 1625	2
	 ("00000000000000000000000000000001"),	 -- 1624	1
	 ("00000000000000000000000000001000"),	 -- 1623	8
	 ("00000000000000000000000000000111"),	 -- 1622	7
	 ("00000000000000000000000000000110"),	 -- 1621	6
	 ("00000000000000000000000000000101"),	 -- 1620	5
	 ("00000000000000000000000000000100"),	 -- 1619	4
	 ("00000000000000000000000000000011"),	 -- 1618	3
	 ("00000000000000000000000000000010"),	 -- 1617	2
	 ("00000000000000000000000000000001"),	 -- 1616	1
	 ("00000000000000000000000000001000"),	 -- 1615	8
	 ("00000000000000000000000000000111"),	 -- 1614	7
	 ("00000000000000000000000000000110"),	 -- 1613	6
	 ("00000000000000000000000000000101"),	 -- 1612	5
	 ("00000000000000000000000000000100"),	 -- 1611	4
	 ("00000000000000000000000000000011"),	 -- 1610	3
	 ("00000000000000000000000000000010"),	 -- 1609	2
	 ("00000000000000000000000000000001"),	 -- 1608	1
	 ("00000000000000000000000000001000"),	 -- 1607	8
	 ("00000000000000000000000000000111"),	 -- 1606	7
	 ("00000000000000000000000000000110"),	 -- 1605	6
	 ("00000000000000000000000000000101"),	 -- 1604	5
	 ("00000000000000000000000000000100"),	 -- 1603	4
	 ("00000000000000000000000000000011"),	 -- 1602	3
	 ("00000000000000000000000000000010"),	 -- 1601	2
	 ("00000000000000000000000000000001"),	 -- 1600	1
	 ("00000000000000000000000000001000"),	 -- 1599	8
	 ("00000000000000000000000000000111"),	 -- 1598	7
	 ("00000000000000000000000000000110"),	 -- 1597	6
	 ("00000000000000000000000000000101"),	 -- 1596	5
	 ("00000000000000000000000000000100"),	 -- 1595	4
	 ("00000000000000000000000000000011"),	 -- 1594	3
	 ("00000000000000000000000000000010"),	 -- 1593	2
	 ("00000000000000000000000000000001"),	 -- 1592	1
	 ("00000000000000000000000000001000"),	 -- 1591	8
	 ("00000000000000000000000000000111"),	 -- 1590	7
	 ("00000000000000000000000000000110"),	 -- 1589	6
	 ("00000000000000000000000000000101"),	 -- 1588	5
	 ("00000000000000000000000000000100"),	 -- 1587	4
	 ("00000000000000000000000000000011"),	 -- 1586	3
	 ("00000000000000000000000000000010"),	 -- 1585	2
	 ("00000000000000000000000000000001"),	 -- 1584	1
	 ("00000000000000000000000000001000"),	 -- 1583	8
	 ("00000000000000000000000000000111"),	 -- 1582	7
	 ("00000000000000000000000000000110"),	 -- 1581	6
	 ("00000000000000000000000000000101"),	 -- 1580	5
	 ("00000000000000000000000000000100"),	 -- 1579	4
	 ("00000000000000000000000000000011"),	 -- 1578	3
	 ("00000000000000000000000000000010"),	 -- 1577	2
	 ("00000000000000000000000000000001"),	 -- 1576	1
	 ("00000000000000000000000000001000"),	 -- 1575	8
	 ("00000000000000000000000000000111"),	 -- 1574	7
	 ("00000000000000000000000000000110"),	 -- 1573	6
	 ("00000000000000000000000000000101"),	 -- 1572	5
	 ("00000000000000000000000000000100"),	 -- 1571	4
	 ("00000000000000000000000000000011"),	 -- 1570	3
	 ("00000000000000000000000000000010"),	 -- 1569	2
	 ("00000000000000000000000000000001"),	 -- 1568	1
	 ("00000000000000000000000000001000"),	 -- 1567	8
	 ("00000000000000000000000000000111"),	 -- 1566	7
	 ("00000000000000000000000000000110"),	 -- 1565	6
	 ("00000000000000000000000000000101"),	 -- 1564	5
	 ("00000000000000000000000000000100"),	 -- 1563	4
	 ("00000000000000000000000000000011"),	 -- 1562	3
	 ("00000000000000000000000000000010"),	 -- 1561	2
	 ("00000000000000000000000000000001"),	 -- 1560	1
	 ("00000000000000000000000000001000"),	 -- 1559	8
	 ("00000000000000000000000000000111"),	 -- 1558	7
	 ("00000000000000000000000000000110"),	 -- 1557	6
	 ("00000000000000000000000000000101"),	 -- 1556	5
	 ("00000000000000000000000000000100"),	 -- 1555	4
	 ("00000000000000000000000000000011"),	 -- 1554	3
	 ("00000000000000000000000000000010"),	 -- 1553	2
	 ("00000000000000000000000000000001"),	 -- 1552	1
	 ("00000000000000000000000000001000"),	 -- 1551	8
	 ("00000000000000000000000000000111"),	 -- 1550	7
	 ("00000000000000000000000000000110"),	 -- 1549	6
	 ("00000000000000000000000000000101"),	 -- 1548	5
	 ("00000000000000000000000000000100"),	 -- 1547	4
	 ("00000000000000000000000000000011"),	 -- 1546	3
	 ("00000000000000000000000000000010"),	 -- 1545	2
	 ("00000000000000000000000000000001"),	 -- 1544	1
	 ("00000000000000000000000000001000"),	 -- 1543	8
	 ("00000000000000000000000000000111"),	 -- 1542	7
	 ("00000000000000000000000000000110"),	 -- 1541	6
	 ("00000000000000000000000000000101"),	 -- 1540	5
	 ("00000000000000000000000000000100"),	 -- 1539	4
	 ("00000000000000000000000000000011"),	 -- 1538	3
	 ("00000000000000000000000000000010"),	 -- 1537	2
	 ("00000000000000000000000000000001"),	 -- 1536	1
	 ("00000000000000000000000000001000"),	 -- 1535	8
	 ("00000000000000000000000000000111"),	 -- 1534	7
	 ("00000000000000000000000000000110"),	 -- 1533	6
	 ("00000000000000000000000000000101"),	 -- 1532	5
	 ("00000000000000000000000000000100"),	 -- 1531	4
	 ("00000000000000000000000000000011"),	 -- 1530	3
	 ("00000000000000000000000000000010"),	 -- 1529	2
	 ("00000000000000000000000000000001"),	 -- 1528	1
	 ("00000000000000000000000000001000"),	 -- 1527	8
	 ("00000000000000000000000000000111"),	 -- 1526	7
	 ("00000000000000000000000000000110"),	 -- 1525	6
	 ("00000000000000000000000000000101"),	 -- 1524	5
	 ("00000000000000000000000000000100"),	 -- 1523	4
	 ("00000000000000000000000000000011"),	 -- 1522	3
	 ("00000000000000000000000000000010"),	 -- 1521	2
	 ("00000000000000000000000000000001"),	 -- 1520	1
	 ("00000000000000000000000000001000"),	 -- 1519	8
	 ("00000000000000000000000000000111"),	 -- 1518	7
	 ("00000000000000000000000000000110"),	 -- 1517	6
	 ("00000000000000000000000000000101"),	 -- 1516	5
	 ("00000000000000000000000000000100"),	 -- 1515	4
	 ("00000000000000000000000000000011"),	 -- 1514	3
	 ("00000000000000000000000000000010"),	 -- 1513	2
	 ("00000000000000000000000000000001"),	 -- 1512	1
	 ("00000000000000000000000000001000"),	 -- 1511	8
	 ("00000000000000000000000000000111"),	 -- 1510	7
	 ("00000000000000000000000000000110"),	 -- 1509	6
	 ("00000000000000000000000000000101"),	 -- 1508	5
	 ("00000000000000000000000000000100"),	 -- 1507	4
	 ("00000000000000000000000000000011"),	 -- 1506	3
	 ("00000000000000000000000000000010"),	 -- 1505	2
	 ("00000000000000000000000000000001"),	 -- 1504	1
	 ("00000000000000000000000000001000"),	 -- 1503	8
	 ("00000000000000000000000000000111"),	 -- 1502	7
	 ("00000000000000000000000000000110"),	 -- 1501	6
	 ("00000000000000000000000000000101"),	 -- 1500	5
	 ("00000000000000000000000000000100"),	 -- 1499	4
	 ("00000000000000000000000000000011"),	 -- 1498	3
	 ("00000000000000000000000000000010"),	 -- 1497	2
	 ("00000000000000000000000000000001"),	 -- 1496	1
	 ("00000000000000000000000000001000"),	 -- 1495	8
	 ("00000000000000000000000000000111"),	 -- 1494	7
	 ("00000000000000000000000000000110"),	 -- 1493	6
	 ("00000000000000000000000000000101"),	 -- 1492	5
	 ("00000000000000000000000000000100"),	 -- 1491	4
	 ("00000000000000000000000000000011"),	 -- 1490	3
	 ("00000000000000000000000000000010"),	 -- 1489	2
	 ("00000000000000000000000000000001"),	 -- 1488	1
	 ("00000000000000000000000000001000"),	 -- 1487	8
	 ("00000000000000000000000000000111"),	 -- 1486	7
	 ("00000000000000000000000000000110"),	 -- 1485	6
	 ("00000000000000000000000000000101"),	 -- 1484	5
	 ("00000000000000000000000000000100"),	 -- 1483	4
	 ("00000000000000000000000000000011"),	 -- 1482	3
	 ("00000000000000000000000000000010"),	 -- 1481	2
	 ("00000000000000000000000000000001"),	 -- 1480	1
	 ("00000000000000000000000000001000"),	 -- 1479	8
	 ("00000000000000000000000000000111"),	 -- 1478	7
	 ("00000000000000000000000000000110"),	 -- 1477	6
	 ("00000000000000000000000000000101"),	 -- 1476	5
	 ("00000000000000000000000000000100"),	 -- 1475	4
	 ("00000000000000000000000000000011"),	 -- 1474	3
	 ("00000000000000000000000000000010"),	 -- 1473	2
	 ("00000000000000000000000000000001"),	 -- 1472	1
	 ("00000000000000000000000000001000"),	 -- 1471	8
	 ("00000000000000000000000000000111"),	 -- 1470	7
	 ("00000000000000000000000000000110"),	 -- 1469	6
	 ("00000000000000000000000000000101"),	 -- 1468	5
	 ("00000000000000000000000000000100"),	 -- 1467	4
	 ("00000000000000000000000000000011"),	 -- 1466	3
	 ("00000000000000000000000000000010"),	 -- 1465	2
	 ("00000000000000000000000000000001"),	 -- 1464	1
	 ("00000000000000000000000000001000"),	 -- 1463	8
	 ("00000000000000000000000000000111"),	 -- 1462	7
	 ("00000000000000000000000000000110"),	 -- 1461	6
	 ("00000000000000000000000000000101"),	 -- 1460	5
	 ("00000000000000000000000000000100"),	 -- 1459	4
	 ("00000000000000000000000000000011"),	 -- 1458	3
	 ("00000000000000000000000000000010"),	 -- 1457	2
	 ("00000000000000000000000000000001"),	 -- 1456	1
	 ("00000000000000000000000000001000"),	 -- 1455	8
	 ("00000000000000000000000000000111"),	 -- 1454	7
	 ("00000000000000000000000000000110"),	 -- 1453	6
	 ("00000000000000000000000000000101"),	 -- 1452	5
	 ("00000000000000000000000000000100"),	 -- 1451	4
	 ("00000000000000000000000000000011"),	 -- 1450	3
	 ("00000000000000000000000000000010"),	 -- 1449	2
	 ("00000000000000000000000000000001"),	 -- 1448	1
	 ("00000000000000000000000000001000"),	 -- 1447	8
	 ("00000000000000000000000000000111"),	 -- 1446	7
	 ("00000000000000000000000000000110"),	 -- 1445	6
	 ("00000000000000000000000000000101"),	 -- 1444	5
	 ("00000000000000000000000000000100"),	 -- 1443	4
	 ("00000000000000000000000000000011"),	 -- 1442	3
	 ("00000000000000000000000000000010"),	 -- 1441	2
	 ("00000000000000000000000000000001"),	 -- 1440	1
	 ("00000000000000000000000000001000"),	 -- 1439	8
	 ("00000000000000000000000000000111"),	 -- 1438	7
	 ("00000000000000000000000000000110"),	 -- 1437	6
	 ("00000000000000000000000000000101"),	 -- 1436	5
	 ("00000000000000000000000000000100"),	 -- 1435	4
	 ("00000000000000000000000000000011"),	 -- 1434	3
	 ("00000000000000000000000000000010"),	 -- 1433	2
	 ("00000000000000000000000000000001"),	 -- 1432	1
	 ("00000000000000000000000000001000"),	 -- 1431	8
	 ("00000000000000000000000000000111"),	 -- 1430	7
	 ("00000000000000000000000000000110"),	 -- 1429	6
	 ("00000000000000000000000000000101"),	 -- 1428	5
	 ("00000000000000000000000000000100"),	 -- 1427	4
	 ("00000000000000000000000000000011"),	 -- 1426	3
	 ("00000000000000000000000000000010"),	 -- 1425	2
	 ("00000000000000000000000000000001"),	 -- 1424	1
	 ("00000000000000000000000000001000"),	 -- 1423	8
	 ("00000000000000000000000000000111"),	 -- 1422	7
	 ("00000000000000000000000000000110"),	 -- 1421	6
	 ("00000000000000000000000000000101"),	 -- 1420	5
	 ("00000000000000000000000000000100"),	 -- 1419	4
	 ("00000000000000000000000000000011"),	 -- 1418	3
	 ("00000000000000000000000000000010"),	 -- 1417	2
	 ("00000000000000000000000000000001"),	 -- 1416	1
	 ("00000000000000000000000000001000"),	 -- 1415	8
	 ("00000000000000000000000000000111"),	 -- 1414	7
	 ("00000000000000000000000000000110"),	 -- 1413	6
	 ("00000000000000000000000000000101"),	 -- 1412	5
	 ("00000000000000000000000000000100"),	 -- 1411	4
	 ("00000000000000000000000000000011"),	 -- 1410	3
	 ("00000000000000000000000000000010"),	 -- 1409	2
	 ("00000000000000000000000000000001"),	 -- 1408	1
	 ("00000000000000000000000000001000"),	 -- 1407	8
	 ("00000000000000000000000000000111"),	 -- 1406	7
	 ("00000000000000000000000000000110"),	 -- 1405	6
	 ("00000000000000000000000000000101"),	 -- 1404	5
	 ("00000000000000000000000000000100"),	 -- 1403	4
	 ("00000000000000000000000000000011"),	 -- 1402	3
	 ("00000000000000000000000000000010"),	 -- 1401	2
	 ("00000000000000000000000000000001"),	 -- 1400	1
	 ("00000000000000000000000000001000"),	 -- 1399	8
	 ("00000000000000000000000000000111"),	 -- 1398	7
	 ("00000000000000000000000000000110"),	 -- 1397	6
	 ("00000000000000000000000000000101"),	 -- 1396	5
	 ("00000000000000000000000000000100"),	 -- 1395	4
	 ("00000000000000000000000000000011"),	 -- 1394	3
	 ("00000000000000000000000000000010"),	 -- 1393	2
	 ("00000000000000000000000000000001"),	 -- 1392	1
	 ("00000000000000000000000000001000"),	 -- 1391	8
	 ("00000000000000000000000000000111"),	 -- 1390	7
	 ("00000000000000000000000000000110"),	 -- 1389	6
	 ("00000000000000000000000000000101"),	 -- 1388	5
	 ("00000000000000000000000000000100"),	 -- 1387	4
	 ("00000000000000000000000000000011"),	 -- 1386	3
	 ("00000000000000000000000000000010"),	 -- 1385	2
	 ("00000000000000000000000000000001"),	 -- 1384	1
	 ("00000000000000000000000000001000"),	 -- 1383	8
	 ("00000000000000000000000000000111"),	 -- 1382	7
	 ("00000000000000000000000000000110"),	 -- 1381	6
	 ("00000000000000000000000000000101"),	 -- 1380	5
	 ("00000000000000000000000000000100"),	 -- 1379	4
	 ("00000000000000000000000000000011"),	 -- 1378	3
	 ("00000000000000000000000000000010"),	 -- 1377	2
	 ("00000000000000000000000000000001"),	 -- 1376	1
	 ("00000000000000000000000000001000"),	 -- 1375	8
	 ("00000000000000000000000000000111"),	 -- 1374	7
	 ("00000000000000000000000000000110"),	 -- 1373	6
	 ("00000000000000000000000000000101"),	 -- 1372	5
	 ("00000000000000000000000000000100"),	 -- 1371	4
	 ("00000000000000000000000000000011"),	 -- 1370	3
	 ("00000000000000000000000000000010"),	 -- 1369	2
	 ("00000000000000000000000000000001"),	 -- 1368	1
	 ("00000000000000000000000000001000"),	 -- 1367	8
	 ("00000000000000000000000000000111"),	 -- 1366	7
	 ("00000000000000000000000000000110"),	 -- 1365	6
	 ("00000000000000000000000000000101"),	 -- 1364	5
	 ("00000000000000000000000000000100"),	 -- 1363	4
	 ("00000000000000000000000000000011"),	 -- 1362	3
	 ("00000000000000000000000000000010"),	 -- 1361	2
	 ("00000000000000000000000000000001"),	 -- 1360	1
	 ("00000000000000000000000000001000"),	 -- 1359	8
	 ("00000000000000000000000000000111"),	 -- 1358	7
	 ("00000000000000000000000000000110"),	 -- 1357	6
	 ("00000000000000000000000000000101"),	 -- 1356	5
	 ("00000000000000000000000000000100"),	 -- 1355	4
	 ("00000000000000000000000000000011"),	 -- 1354	3
	 ("00000000000000000000000000000010"),	 -- 1353	2
	 ("00000000000000000000000000000001"),	 -- 1352	1
	 ("00000000000000000000000000001000"),	 -- 1351	8
	 ("00000000000000000000000000000111"),	 -- 1350	7
	 ("00000000000000000000000000000110"),	 -- 1349	6
	 ("00000000000000000000000000000101"),	 -- 1348	5
	 ("00000000000000000000000000000100"),	 -- 1347	4
	 ("00000000000000000000000000000011"),	 -- 1346	3
	 ("00000000000000000000000000000010"),	 -- 1345	2
	 ("00000000000000000000000000000001"),	 -- 1344	1
	 ("00000000000000000000000000001000"),	 -- 1343	8
	 ("00000000000000000000000000000111"),	 -- 1342	7
	 ("00000000000000000000000000000110"),	 -- 1341	6
	 ("00000000000000000000000000000101"),	 -- 1340	5
	 ("00000000000000000000000000000100"),	 -- 1339	4
	 ("00000000000000000000000000000011"),	 -- 1338	3
	 ("00000000000000000000000000000010"),	 -- 1337	2
	 ("00000000000000000000000000000001"),	 -- 1336	1
	 ("00000000000000000000000000001000"),	 -- 1335	8
	 ("00000000000000000000000000000111"),	 -- 1334	7
	 ("00000000000000000000000000000110"),	 -- 1333	6
	 ("00000000000000000000000000000101"),	 -- 1332	5
	 ("00000000000000000000000000000100"),	 -- 1331	4
	 ("00000000000000000000000000000011"),	 -- 1330	3
	 ("00000000000000000000000000000010"),	 -- 1329	2
	 ("00000000000000000000000000000001"),	 -- 1328	1
	 ("00000000000000000000000000001000"),	 -- 1327	8
	 ("00000000000000000000000000000111"),	 -- 1326	7
	 ("00000000000000000000000000000110"),	 -- 1325	6
	 ("00000000000000000000000000000101"),	 -- 1324	5
	 ("00000000000000000000000000000100"),	 -- 1323	4
	 ("00000000000000000000000000000011"),	 -- 1322	3
	 ("00000000000000000000000000000010"),	 -- 1321	2
	 ("00000000000000000000000000000001"),	 -- 1320	1
	 ("00000000000000000000000000001000"),	 -- 1319	8
	 ("00000000000000000000000000000111"),	 -- 1318	7
	 ("00000000000000000000000000000110"),	 -- 1317	6
	 ("00000000000000000000000000000101"),	 -- 1316	5
	 ("00000000000000000000000000000100"),	 -- 1315	4
	 ("00000000000000000000000000000011"),	 -- 1314	3
	 ("00000000000000000000000000000010"),	 -- 1313	2
	 ("00000000000000000000000000000001"),	 -- 1312	1
	 ("00000000000000000000000000001000"),	 -- 1311	8
	 ("00000000000000000000000000000111"),	 -- 1310	7
	 ("00000000000000000000000000000110"),	 -- 1309	6
	 ("00000000000000000000000000000101"),	 -- 1308	5
	 ("00000000000000000000000000000100"),	 -- 1307	4
	 ("00000000000000000000000000000011"),	 -- 1306	3
	 ("00000000000000000000000000000010"),	 -- 1305	2
	 ("00000000000000000000000000000001"),	 -- 1304	1
	 ("00000000000000000000000000001000"),	 -- 1303	8
	 ("00000000000000000000000000000111"),	 -- 1302	7
	 ("00000000000000000000000000000110"),	 -- 1301	6
	 ("00000000000000000000000000000101"),	 -- 1300	5
	 ("00000000000000000000000000000100"),	 -- 1299	4
	 ("00000000000000000000000000000011"),	 -- 1298	3
	 ("00000000000000000000000000000010"),	 -- 1297	2
	 ("00000000000000000000000000000001"),	 -- 1296	1
	 ("00000000000000000000000000001000"),	 -- 1295	8
	 ("00000000000000000000000000000111"),	 -- 1294	7
	 ("00000000000000000000000000000110"),	 -- 1293	6
	 ("00000000000000000000000000000101"),	 -- 1292	5
	 ("00000000000000000000000000000100"),	 -- 1291	4
	 ("00000000000000000000000000000011"),	 -- 1290	3
	 ("00000000000000000000000000000010"),	 -- 1289	2
	 ("00000000000000000000000000000001"),	 -- 1288	1
	 ("00000000000000000000000000001000"),	 -- 1287	8
	 ("00000000000000000000000000000111"),	 -- 1286	7
	 ("00000000000000000000000000000110"),	 -- 1285	6
	 ("00000000000000000000000000000101"),	 -- 1284	5
	 ("00000000000000000000000000000100"),	 -- 1283	4
	 ("00000000000000000000000000000011"),	 -- 1282	3
	 ("00000000000000000000000000000010"),	 -- 1281	2
	 ("00000000000000000000000000000001"),	 -- 1280	1
	 ("00000000000000000000000000001000"),	 -- 1279	8
	 ("00000000000000000000000000000111"),	 -- 1278	7
	 ("00000000000000000000000000000110"),	 -- 1277	6
	 ("00000000000000000000000000000101"),	 -- 1276	5
	 ("00000000000000000000000000000100"),	 -- 1275	4
	 ("00000000000000000000000000000011"),	 -- 1274	3
	 ("00000000000000000000000000000010"),	 -- 1273	2
	 ("00000000000000000000000000000001"),	 -- 1272	1
	 ("00000000000000000000000000001000"),	 -- 1271	8
	 ("00000000000000000000000000000111"),	 -- 1270	7
	 ("00000000000000000000000000000110"),	 -- 1269	6
	 ("00000000000000000000000000000101"),	 -- 1268	5
	 ("00000000000000000000000000000100"),	 -- 1267	4
	 ("00000000000000000000000000000011"),	 -- 1266	3
	 ("00000000000000000000000000000010"),	 -- 1265	2
	 ("00000000000000000000000000000001"),	 -- 1264	1
	 ("00000000000000000000000000001000"),	 -- 1263	8
	 ("00000000000000000000000000000111"),	 -- 1262	7
	 ("00000000000000000000000000000110"),	 -- 1261	6
	 ("00000000000000000000000000000101"),	 -- 1260	5
	 ("00000000000000000000000000000100"),	 -- 1259	4
	 ("00000000000000000000000000000011"),	 -- 1258	3
	 ("00000000000000000000000000000010"),	 -- 1257	2
	 ("00000000000000000000000000000001"),	 -- 1256	1
	 ("00000000000000000000000000001000"),	 -- 1255	8
	 ("00000000000000000000000000000111"),	 -- 1254	7
	 ("00000000000000000000000000000110"),	 -- 1253	6
	 ("00000000000000000000000000000101"),	 -- 1252	5
	 ("00000000000000000000000000000100"),	 -- 1251	4
	 ("00000000000000000000000000000011"),	 -- 1250	3
	 ("00000000000000000000000000000010"),	 -- 1249	2
	 ("00000000000000000000000000000001"),	 -- 1248	1
	 ("00000000000000000000000000001000"),	 -- 1247	8
	 ("00000000000000000000000000000111"),	 -- 1246	7
	 ("00000000000000000000000000000110"),	 -- 1245	6
	 ("00000000000000000000000000000101"),	 -- 1244	5
	 ("00000000000000000000000000000100"),	 -- 1243	4
	 ("00000000000000000000000000000011"),	 -- 1242	3
	 ("00000000000000000000000000000010"),	 -- 1241	2
	 ("00000000000000000000000000000001"),	 -- 1240	1
	 ("00000000000000000000000000001000"),	 -- 1239	8
	 ("00000000000000000000000000000111"),	 -- 1238	7
	 ("00000000000000000000000000000110"),	 -- 1237	6
	 ("00000000000000000000000000000101"),	 -- 1236	5
	 ("00000000000000000000000000000100"),	 -- 1235	4
	 ("00000000000000000000000000000011"),	 -- 1234	3
	 ("00000000000000000000000000000010"),	 -- 1233	2
	 ("00000000000000000000000000000001"),	 -- 1232	1
	 ("00000000000000000000000000001000"),	 -- 1231	8
	 ("00000000000000000000000000000111"),	 -- 1230	7
	 ("00000000000000000000000000000110"),	 -- 1229	6
	 ("00000000000000000000000000000101"),	 -- 1228	5
	 ("00000000000000000000000000000100"),	 -- 1227	4
	 ("00000000000000000000000000000011"),	 -- 1226	3
	 ("00000000000000000000000000000010"),	 -- 1225	2
	 ("00000000000000000000000000000001"),	 -- 1224	1
	 ("00000000000000000000000000001000"),	 -- 1223	8
	 ("00000000000000000000000000000111"),	 -- 1222	7
	 ("00000000000000000000000000000110"),	 -- 1221	6
	 ("00000000000000000000000000000101"),	 -- 1220	5
	 ("00000000000000000000000000000100"),	 -- 1219	4
	 ("00000000000000000000000000000011"),	 -- 1218	3
	 ("00000000000000000000000000000010"),	 -- 1217	2
	 ("00000000000000000000000000000001"),	 -- 1216	1
	 ("00000000000000000000000000001000"),	 -- 1215	8
	 ("00000000000000000000000000000111"),	 -- 1214	7
	 ("00000000000000000000000000000110"),	 -- 1213	6
	 ("00000000000000000000000000000101"),	 -- 1212	5
	 ("00000000000000000000000000000100"),	 -- 1211	4
	 ("00000000000000000000000000000011"),	 -- 1210	3
	 ("00000000000000000000000000000010"),	 -- 1209	2
	 ("00000000000000000000000000000001"),	 -- 1208	1
	 ("00000000000000000000000000001000"),	 -- 1207	8
	 ("00000000000000000000000000000111"),	 -- 1206	7
	 ("00000000000000000000000000000110"),	 -- 1205	6
	 ("00000000000000000000000000000101"),	 -- 1204	5
	 ("00000000000000000000000000000100"),	 -- 1203	4
	 ("00000000000000000000000000000011"),	 -- 1202	3
	 ("00000000000000000000000000000010"),	 -- 1201	2
	 ("00000000000000000000000000000001"),	 -- 1200	1
	 ("00000000000000000000000000001000"),	 -- 1199	8
	 ("00000000000000000000000000000111"),	 -- 1198	7
	 ("00000000000000000000000000000110"),	 -- 1197	6
	 ("00000000000000000000000000000101"),	 -- 1196	5
	 ("00000000000000000000000000000100"),	 -- 1195	4
	 ("00000000000000000000000000000011"),	 -- 1194	3
	 ("00000000000000000000000000000010"),	 -- 1193	2
	 ("00000000000000000000000000000001"),	 -- 1192	1
	 ("00000000000000000000000000001000"),	 -- 1191	8
	 ("00000000000000000000000000000111"),	 -- 1190	7
	 ("00000000000000000000000000000110"),	 -- 1189	6
	 ("00000000000000000000000000000101"),	 -- 1188	5
	 ("00000000000000000000000000000100"),	 -- 1187	4
	 ("00000000000000000000000000000011"),	 -- 1186	3
	 ("00000000000000000000000000000010"),	 -- 1185	2
	 ("00000000000000000000000000000001"),	 -- 1184	1
	 ("00000000000000000000000000001000"),	 -- 1183	8
	 ("00000000000000000000000000000111"),	 -- 1182	7
	 ("00000000000000000000000000000110"),	 -- 1181	6
	 ("00000000000000000000000000000101"),	 -- 1180	5
	 ("00000000000000000000000000000100"),	 -- 1179	4
	 ("00000000000000000000000000000011"),	 -- 1178	3
	 ("00000000000000000000000000000010"),	 -- 1177	2
	 ("00000000000000000000000000000001"),	 -- 1176	1
	 ("00000000000000000000000000001000"),	 -- 1175	8
	 ("00000000000000000000000000000111"),	 -- 1174	7
	 ("00000000000000000000000000000110"),	 -- 1173	6
	 ("00000000000000000000000000000101"),	 -- 1172	5
	 ("00000000000000000000000000000100"),	 -- 1171	4
	 ("00000000000000000000000000000011"),	 -- 1170	3
	 ("00000000000000000000000000000010"),	 -- 1169	2
	 ("00000000000000000000000000000001"),	 -- 1168	1
	 ("00000000000000000000000000001000"),	 -- 1167	8
	 ("00000000000000000000000000000111"),	 -- 1166	7
	 ("00000000000000000000000000000110"),	 -- 1165	6
	 ("00000000000000000000000000000101"),	 -- 1164	5
	 ("00000000000000000000000000000100"),	 -- 1163	4
	 ("00000000000000000000000000000011"),	 -- 1162	3
	 ("00000000000000000000000000000010"),	 -- 1161	2
	 ("00000000000000000000000000000001"),	 -- 1160	1
	 ("00000000000000000000000000001000"),	 -- 1159	8
	 ("00000000000000000000000000000111"),	 -- 1158	7
	 ("00000000000000000000000000000110"),	 -- 1157	6
	 ("00000000000000000000000000000101"),	 -- 1156	5
	 ("00000000000000000000000000000100"),	 -- 1155	4
	 ("00000000000000000000000000000011"),	 -- 1154	3
	 ("00000000000000000000000000000010"),	 -- 1153	2
	 ("00000000000000000000000000000001"),	 -- 1152	1
	 ("00000000000000000000000000001000"),	 -- 1151	8
	 ("00000000000000000000000000000111"),	 -- 1150	7
	 ("00000000000000000000000000000110"),	 -- 1149	6
	 ("00000000000000000000000000000101"),	 -- 1148	5
	 ("00000000000000000000000000000100"),	 -- 1147	4
	 ("00000000000000000000000000000011"),	 -- 1146	3
	 ("00000000000000000000000000000010"),	 -- 1145	2
	 ("00000000000000000000000000000001"),	 -- 1144	1
	 ("00000000000000000000000000001000"),	 -- 1143	8
	 ("00000000000000000000000000000111"),	 -- 1142	7
	 ("00000000000000000000000000000110"),	 -- 1141	6
	 ("00000000000000000000000000000101"),	 -- 1140	5
	 ("00000000000000000000000000000100"),	 -- 1139	4
	 ("00000000000000000000000000000011"),	 -- 1138	3
	 ("00000000000000000000000000000010"),	 -- 1137	2
	 ("00000000000000000000000000000001"),	 -- 1136	1
	 ("00000000000000000000000000001000"),	 -- 1135	8
	 ("00000000000000000000000000000111"),	 -- 1134	7
	 ("00000000000000000000000000000110"),	 -- 1133	6
	 ("00000000000000000000000000000101"),	 -- 1132	5
	 ("00000000000000000000000000000100"),	 -- 1131	4
	 ("00000000000000000000000000000011"),	 -- 1130	3
	 ("00000000000000000000000000000010"),	 -- 1129	2
	 ("00000000000000000000000000000001"),	 -- 1128	1
	 ("00000000000000000000000000001000"),	 -- 1127	8
	 ("00000000000000000000000000000111"),	 -- 1126	7
	 ("00000000000000000000000000000110"),	 -- 1125	6
	 ("00000000000000000000000000000101"),	 -- 1124	5
	 ("00000000000000000000000000000100"),	 -- 1123	4
	 ("00000000000000000000000000000011"),	 -- 1122	3
	 ("00000000000000000000000000000010"),	 -- 1121	2
	 ("00000000000000000000000000000001"),	 -- 1120	1
	 ("00000000000000000000000000001000"),	 -- 1119	8
	 ("00000000000000000000000000000111"),	 -- 1118	7
	 ("00000000000000000000000000000110"),	 -- 1117	6
	 ("00000000000000000000000000000101"),	 -- 1116	5
	 ("00000000000000000000000000000100"),	 -- 1115	4
	 ("00000000000000000000000000000011"),	 -- 1114	3
	 ("00000000000000000000000000000010"),	 -- 1113	2
	 ("00000000000000000000000000000001"),	 -- 1112	1
	 ("00000000000000000000000000001000"),	 -- 1111	8
	 ("00000000000000000000000000000111"),	 -- 1110	7
	 ("00000000000000000000000000000110"),	 -- 1109	6
	 ("00000000000000000000000000000101"),	 -- 1108	5
	 ("00000000000000000000000000000100"),	 -- 1107	4
	 ("00000000000000000000000000000011"),	 -- 1106	3
	 ("00000000000000000000000000000010"),	 -- 1105	2
	 ("00000000000000000000000000000001"),	 -- 1104	1
	 ("00000000000000000000000000001000"),	 -- 1103	8
	 ("00000000000000000000000000000111"),	 -- 1102	7
	 ("00000000000000000000000000000110"),	 -- 1101	6
	 ("00000000000000000000000000000101"),	 -- 1100	5
	 ("00000000000000000000000000000100"),	 -- 1099	4
	 ("00000000000000000000000000000011"),	 -- 1098	3
	 ("00000000000000000000000000000010"),	 -- 1097	2
	 ("00000000000000000000000000000001"),	 -- 1096	1
	 ("00000000000000000000000000001000"),	 -- 1095	8
	 ("00000000000000000000000000000111"),	 -- 1094	7
	 ("00000000000000000000000000000110"),	 -- 1093	6
	 ("00000000000000000000000000000101"),	 -- 1092	5
	 ("00000000000000000000000000000100"),	 -- 1091	4
	 ("00000000000000000000000000000011"),	 -- 1090	3
	 ("00000000000000000000000000000010"),	 -- 1089	2
	 ("00000000000000000000000000000001"),	 -- 1088	1
	 ("00000000000000000000000000001000"),	 -- 1087	8
	 ("00000000000000000000000000000111"),	 -- 1086	7
	 ("00000000000000000000000000000110"),	 -- 1085	6
	 ("00000000000000000000000000000101"),	 -- 1084	5
	 ("00000000000000000000000000000100"),	 -- 1083	4
	 ("00000000000000000000000000000011"),	 -- 1082	3
	 ("00000000000000000000000000000010"),	 -- 1081	2
	 ("00000000000000000000000000000001"),	 -- 1080	1
	 ("00000000000000000000000000001000"),	 -- 1079	8
	 ("00000000000000000000000000000111"),	 -- 1078	7
	 ("00000000000000000000000000000110"),	 -- 1077	6
	 ("00000000000000000000000000000101"),	 -- 1076	5
	 ("00000000000000000000000000000100"),	 -- 1075	4
	 ("00000000000000000000000000000011"),	 -- 1074	3
	 ("00000000000000000000000000000010"),	 -- 1073	2
	 ("00000000000000000000000000000001"),	 -- 1072	1
	 ("00000000000000000000000000001000"),	 -- 1071	8
	 ("00000000000000000000000000000111"),	 -- 1070	7
	 ("00000000000000000000000000000110"),	 -- 1069	6
	 ("00000000000000000000000000000101"),	 -- 1068	5
	 ("00000000000000000000000000000100"),	 -- 1067	4
	 ("00000000000000000000000000000011"),	 -- 1066	3
	 ("00000000000000000000000000000010"),	 -- 1065	2
	 ("00000000000000000000000000000001"),	 -- 1064	1
	 ("00000000000000000000000000001000"),	 -- 1063	8
	 ("00000000000000000000000000000111"),	 -- 1062	7
	 ("00000000000000000000000000000110"),	 -- 1061	6
	 ("00000000000000000000000000000101"),	 -- 1060	5
	 ("00000000000000000000000000000100"),	 -- 1059	4
	 ("00000000000000000000000000000011"),	 -- 1058	3
	 ("00000000000000000000000000000010"),	 -- 1057	2
	 ("00000000000000000000000000000001"),	 -- 1056	1
	 ("00000000000000000000000000001000"),	 -- 1055	8
	 ("00000000000000000000000000000111"),	 -- 1054	7
	 ("00000000000000000000000000000110"),	 -- 1053	6
	 ("00000000000000000000000000000101"),	 -- 1052	5
	 ("00000000000000000000000000000100"),	 -- 1051	4
	 ("00000000000000000000000000000011"),	 -- 1050	3
	 ("00000000000000000000000000000010"),	 -- 1049	2
	 ("00000000000000000000000000000001"),	 -- 1048	1
	 ("00000000000000000000000000001000"),	 -- 1047	8
	 ("00000000000000000000000000000111"),	 -- 1046	7
	 ("00000000000000000000000000000110"),	 -- 1045	6
	 ("00000000000000000000000000000101"),	 -- 1044	5
	 ("00000000000000000000000000000100"),	 -- 1043	4
	 ("00000000000000000000000000000011"),	 -- 1042	3
	 ("00000000000000000000000000000010"),	 -- 1041	2
	 ("00000000000000000000000000000001"),	 -- 1040	1
	 ("00000000000000000000000000001000"),	 -- 1039	8
	 ("00000000000000000000000000000111"),	 -- 1038	7
	 ("00000000000000000000000000000110"),	 -- 1037	6
	 ("00000000000000000000000000000101"),	 -- 1036	5
	 ("00000000000000000000000000000100"),	 -- 1035	4
	 ("00000000000000000000000000000011"),	 -- 1034	3
	 ("00000000000000000000000000000010"),	 -- 1033	2
	 ("00000000000000000000000000000001"),	 -- 1032	1
	 ("00000000000000000000000000001000"),	 -- 1031	8
	 ("00000000000000000000000000000111"),	 -- 1030	7
	 ("00000000000000000000000000000110"),	 -- 1029	6
	 ("00000000000000000000000000000101"),	 -- 1028	5
	 ("00000000000000000000000000000100"),	 -- 1027	4
	 ("00000000000000000000000000000011"),	 -- 1026	3
	 ("00000000000000000000000000000010"),	 -- 1025	2
	 ("00000000000000000000000000000001"),	 -- 1024	1
	 ("00000000000000000000000001010000"),	 -- 1023	80
	 ("00000000000000000000000000000111"),	 -- 1022	7
	 ("00000000000000000000000000000110"),	 -- 1021	6
	 ("00000000000000000000000000000101"),	 -- 1020	5
	 ("00000000000000000000000000000100"),	 -- 1019	4
	 ("00000000000000000000000000000011"),	 -- 1018	3
	 ("00000000000000000000000000000010"),	 -- 1017	2
	 ("00000000000000000000000000000001"),	 -- 1016	1
	 ("00000000000000000000000000001000"),	 -- 1015	8
	 ("00000000000000000000000000000111"),	 -- 1014	7
	 ("00000000000000000000000000000110"),	 -- 1013	6
	 ("00000000000000000000000000000101"),	 -- 1012	5
	 ("00000000000000000000000000000100"),	 -- 1011	4
	 ("00000000000000000000000000000011"),	 -- 1010	3
	 ("00000000000000000000000000000010"),	 -- 1009	2
	 ("00000000000000000000000000000001"),	 -- 1008	1
	 ("00000000000000000000000000001000"),	 -- 1007	8
	 ("00000000000000000000000000000111"),	 -- 1006	7
	 ("00000000000000000000000000000110"),	 -- 1005	6
	 ("00000000000000000000000000000101"),	 -- 1004	5
	 ("00000000000000000000000000000100"),	 -- 1003	4
	 ("00000000000000000000000000000011"),	 -- 1002	3
	 ("00000000000000000000000000000010"),	 -- 1001	2
	 ("00000000000000000000000000000001"),	 -- 1000	1
	 ("00000000000000000000000000001000"),	 -- 999	8
	 ("00000000000000000000000000000111"),	 -- 998	7
	 ("00000000000000000000000000000110"),	 -- 997	6
	 ("00000000000000000000000000000101"),	 -- 996	5
	 ("00000000000000000000000000000100"),	 -- 995	4
	 ("00000000000000000000000000000011"),	 -- 994	3
	 ("00000000000000000000000000000010"),	 -- 993	2
	 ("00000000000000000000000000000001"),	 -- 992	1
	 ("00000000000000000000000000001000"),	 -- 991	8
	 ("00000000000000000000000000000111"),	 -- 990	7
	 ("00000000000000000000000000000110"),	 -- 989	6
	 ("00000000000000000000000000000101"),	 -- 988	5
	 ("00000000000000000000000000000100"),	 -- 987	4
	 ("00000000000000000000000000000011"),	 -- 986	3
	 ("00000000000000000000000000000010"),	 -- 985	2
	 ("00000000000000000000000000000001"),	 -- 984	1
	 ("00000000000000000000000000001000"),	 -- 983	8
	 ("00000000000000000000000000000111"),	 -- 982	7
	 ("00000000000000000000000000000110"),	 -- 981	6
	 ("00000000000000000000000000000101"),	 -- 980	5
	 ("00000000000000000000000000000100"),	 -- 979	4
	 ("00000000000000000000000000000011"),	 -- 978	3
	 ("00000000000000000000000000000010"),	 -- 977	2
	 ("00000000000000000000000000000001"),	 -- 976	1
	 ("00000000000000000000000000001000"),	 -- 975	8
	 ("00000000000000000000000000000111"),	 -- 974	7
	 ("00000000000000000000000000000110"),	 -- 973	6
	 ("00000000000000000000000000000101"),	 -- 972	5
	 ("00000000000000000000000000000100"),	 -- 971	4
	 ("00000000000000000000000000000011"),	 -- 970	3
	 ("00000000000000000000000000000010"),	 -- 969	2
	 ("00000000000000000000000000000001"),	 -- 968	1
	 ("00000000000000000000000000001000"),	 -- 967	8
	 ("00000000000000000000000000000111"),	 -- 966	7
	 ("00000000000000000000000000000110"),	 -- 965	6
	 ("00000000000000000000000000000101"),	 -- 964	5
	 ("00000000000000000000000000000100"),	 -- 963	4
	 ("00000000000000000000000000000011"),	 -- 962	3
	 ("00000000000000000000000000000010"),	 -- 961	2
	 ("00000000000000000000000000000001"),	 -- 960	1
	 ("00000000000000000000000000001000"),	 -- 959	8
	 ("00000000000000000000000000000111"),	 -- 958	7
	 ("00000000000000000000000000000110"),	 -- 957	6
	 ("00000000000000000000000000000101"),	 -- 956	5
	 ("00000000000000000000000000000100"),	 -- 955	4
	 ("00000000000000000000000000000011"),	 -- 954	3
	 ("00000000000000000000000000000010"),	 -- 953	2
	 ("00000000000000000000000000000001"),	 -- 952	1
	 ("00000000000000000000000000001000"),	 -- 951	8
	 ("00000000000000000000000000000111"),	 -- 950	7
	 ("00000000000000000000000000000110"),	 -- 949	6
	 ("00000000000000000000000000000101"),	 -- 948	5
	 ("00000000000000000000000000000100"),	 -- 947	4
	 ("00000000000000000000000000000011"),	 -- 946	3
	 ("00000000000000000000000000000010"),	 -- 945	2
	 ("00000000000000000000000000000001"),	 -- 944	1
	 ("00000000000000000000000000001000"),	 -- 943	8
	 ("00000000000000000000000000000111"),	 -- 942	7
	 ("00000000000000000000000000000110"),	 -- 941	6
	 ("00000000000000000000000000000101"),	 -- 940	5
	 ("00000000000000000000000000000100"),	 -- 939	4
	 ("00000000000000000000000000000011"),	 -- 938	3
	 ("00000000000000000000000000000010"),	 -- 937	2
	 ("00000000000000000000000000000001"),	 -- 936	1
	 ("00000000000000000000000000001000"),	 -- 935	8
	 ("00000000000000000000000000000111"),	 -- 934	7
	 ("00000000000000000000000000000110"),	 -- 933	6
	 ("00000000000000000000000000000101"),	 -- 932	5
	 ("00000000000000000000000000000100"),	 -- 931	4
	 ("00000000000000000000000000000011"),	 -- 930	3
	 ("00000000000000000000000000000010"),	 -- 929	2
	 ("00000000000000000000000000000001"),	 -- 928	1
	 ("00000000000000000000000000001000"),	 -- 927	8
	 ("00000000000000000000000000000111"),	 -- 926	7
	 ("00000000000000000000000000000110"),	 -- 925	6
	 ("00000000000000000000000000000101"),	 -- 924	5
	 ("00000000000000000000000000000100"),	 -- 923	4
	 ("00000000000000000000000000000011"),	 -- 922	3
	 ("00000000000000000000000000000010"),	 -- 921	2
	 ("00000000000000000000000000000001"),	 -- 920	1
	 ("00000000000000000000000000001000"),	 -- 919	8
	 ("00000000000000000000000000000111"),	 -- 918	7
	 ("00000000000000000000000000000110"),	 -- 917	6
	 ("00000000000000000000000000000101"),	 -- 916	5
	 ("00000000000000000000000000000100"),	 -- 915	4
	 ("00000000000000000000000000000011"),	 -- 914	3
	 ("00000000000000000000000000000010"),	 -- 913	2
	 ("00000000000000000000000000000001"),	 -- 912	1
	 ("00000000000000000000000000001000"),	 -- 911	8
	 ("00000000000000000000000000000111"),	 -- 910	7
	 ("00000000000000000000000000000110"),	 -- 909	6
	 ("00000000000000000000000000000101"),	 -- 908	5
	 ("00000000000000000000000000000100"),	 -- 907	4
	 ("00000000000000000000000000000011"),	 -- 906	3
	 ("00000000000000000000000000000010"),	 -- 905	2
	 ("00000000000000000000000000000001"),	 -- 904	1
	 ("00000000000000000000000000001000"),	 -- 903	8
	 ("00000000000000000000000000000111"),	 -- 902	7
	 ("00000000000000000000000000000110"),	 -- 901	6
	 ("00000000000000000000000000000101"),	 -- 900	5
	 ("00000000000000000000000000000100"),	 -- 899	4
	 ("00000000000000000000000000000011"),	 -- 898	3
	 ("00000000000000000000000000000010"),	 -- 897	2
	 ("00000000000000000000000000000001"),	 -- 896	1
	 ("00000000000000000000000000001000"),	 -- 895	8
	 ("00000000000000000000000000000111"),	 -- 894	7
	 ("00000000000000000000000000000110"),	 -- 893	6
	 ("00000000000000000000000000000101"),	 -- 892	5
	 ("00000000000000000000000000000100"),	 -- 891	4
	 ("00000000000000000000000000000011"),	 -- 890	3
	 ("00000000000000000000000000000010"),	 -- 889	2
	 ("00000000000000000000000000000001"),	 -- 888	1
	 ("00000000000000000000000000001000"),	 -- 887	8
	 ("00000000000000000000000000000111"),	 -- 886	7
	 ("00000000000000000000000000000110"),	 -- 885	6
	 ("00000000000000000000000000000101"),	 -- 884	5
	 ("00000000000000000000000000000100"),	 -- 883	4
	 ("00000000000000000000000000000011"),	 -- 882	3
	 ("00000000000000000000000000000010"),	 -- 881	2
	 ("00000000000000000000000000000001"),	 -- 880	1
	 ("00000000000000000000000000001000"),	 -- 879	8
	 ("00000000000000000000000000000111"),	 -- 878	7
	 ("00000000000000000000000000000110"),	 -- 877	6
	 ("00000000000000000000000000000101"),	 -- 876	5
	 ("00000000000000000000000000000100"),	 -- 875	4
	 ("00000000000000000000000000000011"),	 -- 874	3
	 ("00000000000000000000000000000010"),	 -- 873	2
	 ("00000000000000000000000000000001"),	 -- 872	1
	 ("00000000000000000000000000001000"),	 -- 871	8
	 ("00000000000000000000000000000111"),	 -- 870	7
	 ("00000000000000000000000000000110"),	 -- 869	6
	 ("00000000000000000000000000000101"),	 -- 868	5
	 ("00000000000000000000000000000100"),	 -- 867	4
	 ("00000000000000000000000000000011"),	 -- 866	3
	 ("00000000000000000000000000000010"),	 -- 865	2
	 ("00000000000000000000000000000001"),	 -- 864	1
	 ("00000000000000000000000000001000"),	 -- 863	8
	 ("00000000000000000000000000000111"),	 -- 862	7
	 ("00000000000000000000000000000110"),	 -- 861	6
	 ("00000000000000000000000000000101"),	 -- 860	5
	 ("00000000000000000000000000000100"),	 -- 859	4
	 ("00000000000000000000000000000011"),	 -- 858	3
	 ("00000000000000000000000000000010"),	 -- 857	2
	 ("00000000000000000000000000000001"),	 -- 856	1
	 ("00000000000000000000000000001000"),	 -- 855	8
	 ("00000000000000000000000000000111"),	 -- 854	7
	 ("00000000000000000000000000000110"),	 -- 853	6
	 ("00000000000000000000000000000101"),	 -- 852	5
	 ("00000000000000000000000000000100"),	 -- 851	4
	 ("00000000000000000000000000000011"),	 -- 850	3
	 ("00000000000000000000000000000010"),	 -- 849	2
	 ("00000000000000000000000000000001"),	 -- 848	1
	 ("00000000000000000000000000001000"),	 -- 847	8
	 ("00000000000000000000000000000111"),	 -- 846	7
	 ("00000000000000000000000000000110"),	 -- 845	6
	 ("00000000000000000000000000000101"),	 -- 844	5
	 ("00000000000000000000000000000100"),	 -- 843	4
	 ("00000000000000000000000000000011"),	 -- 842	3
	 ("00000000000000000000000000000010"),	 -- 841	2
	 ("00000000000000000000000000000001"),	 -- 840	1
	 ("00000000000000000000000000001000"),	 -- 839	8
	 ("00000000000000000000000000000111"),	 -- 838	7
	 ("00000000000000000000000000000110"),	 -- 837	6
	 ("00000000000000000000000000000101"),	 -- 836	5
	 ("00000000000000000000000000000100"),	 -- 835	4
	 ("00000000000000000000000000000011"),	 -- 834	3
	 ("00000000000000000000000000000010"),	 -- 833	2
	 ("00000000000000000000000000000001"),	 -- 832	1
	 ("00000000000000000000000000001000"),	 -- 831	8
	 ("00000000000000000000000000000111"),	 -- 830	7
	 ("00000000000000000000000000000110"),	 -- 829	6
	 ("00000000000000000000000000000101"),	 -- 828	5
	 ("00000000000000000000000000000100"),	 -- 827	4
	 ("00000000000000000000000000000011"),	 -- 826	3
	 ("00000000000000000000000000000010"),	 -- 825	2
	 ("00000000000000000000000000000001"),	 -- 824	1
	 ("00000000000000000000000000001000"),	 -- 823	8
	 ("00000000000000000000000000000111"),	 -- 822	7
	 ("00000000000000000000000000000110"),	 -- 821	6
	 ("00000000000000000000000000000101"),	 -- 820	5
	 ("00000000000000000000000000000100"),	 -- 819	4
	 ("00000000000000000000000000000011"),	 -- 818	3
	 ("00000000000000000000000000000010"),	 -- 817	2
	 ("00000000000000000000000000000001"),	 -- 816	1
	 ("00000000000000000000000000001000"),	 -- 815	8
	 ("00000000000000000000000000000111"),	 -- 814	7
	 ("00000000000000000000000000000110"),	 -- 813	6
	 ("00000000000000000000000000000101"),	 -- 812	5
	 ("00000000000000000000000000000100"),	 -- 811	4
	 ("00000000000000000000000000000011"),	 -- 810	3
	 ("00000000000000000000000000000010"),	 -- 809	2
	 ("00000000000000000000000000000001"),	 -- 808	1
	 ("00000000000000000000000000001000"),	 -- 807	8
	 ("00000000000000000000000000000111"),	 -- 806	7
	 ("00000000000000000000000000000110"),	 -- 805	6
	 ("00000000000000000000000000000101"),	 -- 804	5
	 ("00000000000000000000000000000100"),	 -- 803	4
	 ("00000000000000000000000000000011"),	 -- 802	3
	 ("00000000000000000000000000000010"),	 -- 801	2
	 ("00000000000000000000000000000001"),	 -- 800	1
	 ("00000000000000000000000000001000"),	 -- 799	8
	 ("00000000000000000000000000000111"),	 -- 798	7
	 ("00000000000000000000000000000110"),	 -- 797	6
	 ("00000000000000000000000000000101"),	 -- 796	5
	 ("00000000000000000000000000000100"),	 -- 795	4
	 ("00000000000000000000000000000011"),	 -- 794	3
	 ("00000000000000000000000000000010"),	 -- 793	2
	 ("00000000000000000000000000000001"),	 -- 792	1
	 ("00000000000000000000000000001000"),	 -- 791	8
	 ("00000000000000000000000000000111"),	 -- 790	7
	 ("00000000000000000000000000000110"),	 -- 789	6
	 ("00000000000000000000000000000101"),	 -- 788	5
	 ("00000000000000000000000000000100"),	 -- 787	4
	 ("00000000000000000000000000000011"),	 -- 786	3
	 ("00000000000000000000000000000010"),	 -- 785	2
	 ("00000000000000000000000000000001"),	 -- 784	1
	 ("00000000000000000000000000001000"),	 -- 783	8
	 ("00000000000000000000000000000111"),	 -- 782	7
	 ("00000000000000000000000000000110"),	 -- 781	6
	 ("00000000000000000000000000000101"),	 -- 780	5
	 ("00000000000000000000000000000100"),	 -- 779	4
	 ("00000000000000000000000000000011"),	 -- 778	3
	 ("00000000000000000000000000000010"),	 -- 777	2
	 ("00000000000000000000000000000001"),	 -- 776	1
	 ("00000000000000000000000000001000"),	 -- 775	8
	 ("00000000000000000000000000000111"),	 -- 774	7
	 ("00000000000000000000000000000110"),	 -- 773	6
	 ("00000000000000000000000000000101"),	 -- 772	5
	 ("00000000000000000000000000000100"),	 -- 771	4
	 ("00000000000000000000000000000011"),	 -- 770	3
	 ("00000000000000000000000000000010"),	 -- 769	2
	 ("00000000000000000000000000000001"),	 -- 768	1
	 ("00000000000000000000000000001000"),	 -- 767	8
	 ("00000000000000000000000000000111"),	 -- 766	7
	 ("00000000000000000000000000000110"),	 -- 765	6
	 ("00000000000000000000000000000101"),	 -- 764	5
	 ("00000000000000000000000000000100"),	 -- 763	4
	 ("00000000000000000000000000000011"),	 -- 762	3
	 ("00000000000000000000000000000010"),	 -- 761	2
	 ("00000000000000000000000000000001"),	 -- 760	1
	 ("00000000000000000000000000001000"),	 -- 759	8
	 ("00000000000000000000000000000111"),	 -- 758	7
	 ("00000000000000000000000000000110"),	 -- 757	6
	 ("00000000000000000000000000000101"),	 -- 756	5
	 ("00000000000000000000000000000100"),	 -- 755	4
	 ("00000000000000000000000000000011"),	 -- 754	3
	 ("00000000000000000000000000000010"),	 -- 753	2
	 ("00000000000000000000000000000001"),	 -- 752	1
	 ("00000000000000000000000000001000"),	 -- 751	8
	 ("00000000000000000000000000000111"),	 -- 750	7
	 ("00000000000000000000000000000110"),	 -- 749	6
	 ("00000000000000000000000000000101"),	 -- 748	5
	 ("00000000000000000000000000000100"),	 -- 747	4
	 ("00000000000000000000000000000011"),	 -- 746	3
	 ("00000000000000000000000000000010"),	 -- 745	2
	 ("00000000000000000000000000000001"),	 -- 744	1
	 ("00000000000000000000000000001000"),	 -- 743	8
	 ("00000000000000000000000000000111"),	 -- 742	7
	 ("00000000000000000000000000000110"),	 -- 741	6
	 ("00000000000000000000000000000101"),	 -- 740	5
	 ("00000000000000000000000000000100"),	 -- 739	4
	 ("00000000000000000000000000000011"),	 -- 738	3
	 ("00000000000000000000000000000010"),	 -- 737	2
	 ("00000000000000000000000000000001"),	 -- 736	1
	 ("00000000000000000000000000001000"),	 -- 735	8
	 ("00000000000000000000000000000111"),	 -- 734	7
	 ("00000000000000000000000000000110"),	 -- 733	6
	 ("00000000000000000000000000000101"),	 -- 732	5
	 ("00000000000000000000000000000100"),	 -- 731	4
	 ("00000000000000000000000000000011"),	 -- 730	3
	 ("00000000000000000000000000000010"),	 -- 729	2
	 ("00000000000000000000000000000001"),	 -- 728	1
	 ("00000000000000000000000000001000"),	 -- 727	8
	 ("00000000000000000000000000000111"),	 -- 726	7
	 ("00000000000000000000000000000110"),	 -- 725	6
	 ("00000000000000000000000000000101"),	 -- 724	5
	 ("00000000000000000000000000000100"),	 -- 723	4
	 ("00000000000000000000000000000011"),	 -- 722	3
	 ("00000000000000000000000000000010"),	 -- 721	2
	 ("00000000000000000000000000000001"),	 -- 720	1
	 ("00000000000000000000000000001000"),	 -- 719	8
	 ("00000000000000000000000000000111"),	 -- 718	7
	 ("00000000000000000000000000000110"),	 -- 717	6
	 ("00000000000000000000000000000101"),	 -- 716	5
	 ("00000000000000000000000000000100"),	 -- 715	4
	 ("00000000000000000000000000000011"),	 -- 714	3
	 ("00000000000000000000000000000010"),	 -- 713	2
	 ("00000000000000000000000000000001"),	 -- 712	1
	 ("00000000000000000000000000001000"),	 -- 711	8
	 ("00000000000000000000000000000111"),	 -- 710	7
	 ("00000000000000000000000000000110"),	 -- 709	6
	 ("00000000000000000000000000000101"),	 -- 708	5
	 ("00000000000000000000000000000100"),	 -- 707	4
	 ("00000000000000000000000000000011"),	 -- 706	3
	 ("00000000000000000000000000000010"),	 -- 705	2
	 ("00000000000000000000000000000001"),	 -- 704	1
	 ("00000000000000000000000000001000"),	 -- 703	8
	 ("00000000000000000000000000000111"),	 -- 702	7
	 ("00000000000000000000000000000110"),	 -- 701	6
	 ("00000000000000000000000000000101"),	 -- 700	5
	 ("00000000000000000000000000000100"),	 -- 699	4
	 ("00000000000000000000000000000011"),	 -- 698	3
	 ("00000000000000000000000000000010"),	 -- 697	2
	 ("00000000000000000000000000000001"),	 -- 696	1
	 ("00000000000000000000000000001000"),	 -- 695	8
	 ("00000000000000000000000000000111"),	 -- 694	7
	 ("00000000000000000000000000000110"),	 -- 693	6
	 ("00000000000000000000000000000101"),	 -- 692	5
	 ("00000000000000000000000000000100"),	 -- 691	4
	 ("00000000000000000000000000000011"),	 -- 690	3
	 ("00000000000000000000000000000010"),	 -- 689	2
	 ("00000000000000000000000000000001"),	 -- 688	1
	 ("00000000000000000000000000001000"),	 -- 687	8
	 ("00000000000000000000000000000111"),	 -- 686	7
	 ("00000000000000000000000000000110"),	 -- 685	6
	 ("00000000000000000000000000000101"),	 -- 684	5
	 ("00000000000000000000000000000100"),	 -- 683	4
	 ("00000000000000000000000000000011"),	 -- 682	3
	 ("00000000000000000000000000000010"),	 -- 681	2
	 ("00000000000000000000000000000001"),	 -- 680	1
	 ("00000000000000000000000000001000"),	 -- 679	8
	 ("00000000000000000000000000000111"),	 -- 678	7
	 ("00000000000000000000000000000110"),	 -- 677	6
	 ("00000000000000000000000000000101"),	 -- 676	5
	 ("00000000000000000000000000000100"),	 -- 675	4
	 ("00000000000000000000000000000011"),	 -- 674	3
	 ("00000000000000000000000000000010"),	 -- 673	2
	 ("00000000000000000000000000000001"),	 -- 672	1
	 ("00000000000000000000000000001000"),	 -- 671	8
	 ("00000000000000000000000000000111"),	 -- 670	7
	 ("00000000000000000000000000000110"),	 -- 669	6
	 ("00000000000000000000000000000101"),	 -- 668	5
	 ("00000000000000000000000000000100"),	 -- 667	4
	 ("00000000000000000000000000000011"),	 -- 666	3
	 ("00000000000000000000000000000010"),	 -- 665	2
	 ("00000000000000000000000000000001"),	 -- 664	1
	 ("00000000000000000000000000001000"),	 -- 663	8
	 ("00000000000000000000000000000111"),	 -- 662	7
	 ("00000000000000000000000000000110"),	 -- 661	6
	 ("00000000000000000000000000000101"),	 -- 660	5
	 ("00000000000000000000000000000100"),	 -- 659	4
	 ("00000000000000000000000000000011"),	 -- 658	3
	 ("00000000000000000000000000000010"),	 -- 657	2
	 ("00000000000000000000000000000001"),	 -- 656	1
	 ("00000000000000000000000000001000"),	 -- 655	8
	 ("00000000000000000000000000000111"),	 -- 654	7
	 ("00000000000000000000000000000110"),	 -- 653	6
	 ("00000000000000000000000000000101"),	 -- 652	5
	 ("00000000000000000000000000000100"),	 -- 651	4
	 ("00000000000000000000000000000011"),	 -- 650	3
	 ("00000000000000000000000000000010"),	 -- 649	2
	 ("00000000000000000000000000000001"),	 -- 648	1
	 ("00000000000000000000000000001000"),	 -- 647	8
	 ("00000000000000000000000000000111"),	 -- 646	7
	 ("00000000000000000000000000000110"),	 -- 645	6
	 ("00000000000000000000000000000101"),	 -- 644	5
	 ("00000000000000000000000000000100"),	 -- 643	4
	 ("00000000000000000000000000000011"),	 -- 642	3
	 ("00000000000000000000000000000010"),	 -- 641	2
	 ("00000000000000000000000000000001"),	 -- 640	1
	 ("00000000000000000000000000001000"),	 -- 639	8
	 ("00000000000000000000000000000111"),	 -- 638	7
	 ("00000000000000000000000000000110"),	 -- 637	6
	 ("00000000000000000000000000000101"),	 -- 636	5
	 ("00000000000000000000000000000100"),	 -- 635	4
	 ("00000000000000000000000000000011"),	 -- 634	3
	 ("00000000000000000000000000000010"),	 -- 633	2
	 ("00000000000000000000000000000001"),	 -- 632	1
	 ("00000000000000000000000000001000"),	 -- 631	8
	 ("00000000000000000000000000000111"),	 -- 630	7
	 ("00000000000000000000000000000110"),	 -- 629	6
	 ("00000000000000000000000000000101"),	 -- 628	5
	 ("00000000000000000000000000000100"),	 -- 627	4
	 ("00000000000000000000000000000011"),	 -- 626	3
	 ("00000000000000000000000000000010"),	 -- 625	2
	 ("00000000000000000000000000000001"),	 -- 624	1
	 ("00000000000000000000000000001000"),	 -- 623	8
	 ("00000000000000000000000000000111"),	 -- 622	7
	 ("00000000000000000000000000000110"),	 -- 621	6
	 ("00000000000000000000000000000101"),	 -- 620	5
	 ("00000000000000000000000000000100"),	 -- 619	4
	 ("00000000000000000000000000000011"),	 -- 618	3
	 ("00000000000000000000000000000010"),	 -- 617	2
	 ("00000000000000000000000000000001"),	 -- 616	1
	 ("00000000000000000000000000001000"),	 -- 615	8
	 ("00000000000000000000000000000111"),	 -- 614	7
	 ("00000000000000000000000000000110"),	 -- 613	6
	 ("00000000000000000000000000000101"),	 -- 612	5
	 ("00000000000000000000000000000100"),	 -- 611	4
	 ("00000000000000000000000000000011"),	 -- 610	3
	 ("00000000000000000000000000000010"),	 -- 609	2
	 ("00000000000000000000000000000001"),	 -- 608	1
	 ("00000000000000000000000000001000"),	 -- 607	8
	 ("00000000000000000000000000000111"),	 -- 606	7
	 ("00000000000000000000000000000110"),	 -- 605	6
	 ("00000000000000000000000000000101"),	 -- 604	5
	 ("00000000000000000000000000000100"),	 -- 603	4
	 ("00000000000000000000000000000011"),	 -- 602	3
	 ("00000000000000000000000000000010"),	 -- 601	2
	 ("00000000000000000000000000000001"),	 -- 600	1
	 ("00000000000000000000000000001000"),	 -- 599	8
	 ("00000000000000000000000000000111"),	 -- 598	7
	 ("00000000000000000000000000000110"),	 -- 597	6
	 ("00000000000000000000000000000101"),	 -- 596	5
	 ("00000000000000000000000000000100"),	 -- 595	4
	 ("00000000000000000000000000000011"),	 -- 594	3
	 ("00000000000000000000000000000010"),	 -- 593	2
	 ("00000000000000000000000000000001"),	 -- 592	1
	 ("00000000000000000000000000001000"),	 -- 591	8
	 ("00000000000000000000000000000111"),	 -- 590	7
	 ("00000000000000000000000000000110"),	 -- 589	6
	 ("00000000000000000000000000000101"),	 -- 588	5
	 ("00000000000000000000000000000100"),	 -- 587	4
	 ("00000000000000000000000000000011"),	 -- 586	3
	 ("00000000000000000000000000000010"),	 -- 585	2
	 ("00000000000000000000000000000001"),	 -- 584	1
	 ("00000000000000000000000000001000"),	 -- 583	8
	 ("00000000000000000000000000000111"),	 -- 582	7
	 ("00000000000000000000000000000110"),	 -- 581	6
	 ("00000000000000000000000000000101"),	 -- 580	5
	 ("00000000000000000000000000000100"),	 -- 579	4
	 ("00000000000000000000000000000011"),	 -- 578	3
	 ("00000000000000000000000000000010"),	 -- 577	2
	 ("00000000000000000000000000000001"),	 -- 576	1
	 ("00000000000000000000000000001000"),	 -- 575	8
	 ("00000000000000000000000000000111"),	 -- 574	7
	 ("00000000000000000000000000000110"),	 -- 573	6
	 ("00000000000000000000000000000101"),	 -- 572	5
	 ("00000000000000000000000000000100"),	 -- 571	4
	 ("00000000000000000000000000000011"),	 -- 570	3
	 ("00000000000000000000000000000010"),	 -- 569	2
	 ("00000000000000000000000000000001"),	 -- 568	1
	 ("00000000000000000000000000001000"),	 -- 567	8
	 ("00000000000000000000000000000111"),	 -- 566	7
	 ("00000000000000000000000000000110"),	 -- 565	6
	 ("00000000000000000000000000000101"),	 -- 564	5
	 ("00000000000000000000000000000100"),	 -- 563	4
	 ("00000000000000000000000000000011"),	 -- 562	3
	 ("00000000000000000000000000000010"),	 -- 561	2
	 ("00000000000000000000000000000001"),	 -- 560	1
	 ("00000000000000000000000000001000"),	 -- 559	8
	 ("00000000000000000000000000000111"),	 -- 558	7
	 ("00000000000000000000000000000110"),	 -- 557	6
	 ("00000000000000000000000000000101"),	 -- 556	5
	 ("00000000000000000000000000000100"),	 -- 555	4
	 ("00000000000000000000000000000011"),	 -- 554	3
	 ("00000000000000000000000000000010"),	 -- 553	2
	 ("00000000000000000000000000000001"),	 -- 552	1
	 ("00000000000000000000000000001000"),	 -- 551	8
	 ("00000000000000000000000000000111"),	 -- 550	7
	 ("00000000000000000000000000000110"),	 -- 549	6
	 ("00000000000000000000000000000101"),	 -- 548	5
	 ("00000000000000000000000000000100"),	 -- 547	4
	 ("00000000000000000000000000000011"),	 -- 546	3
	 ("00000000000000000000000000000010"),	 -- 545	2
	 ("00000000000000000000000000000001"),	 -- 544	1
	 ("00000000000000000000000000001000"),	 -- 543	8
	 ("00000000000000000000000000000111"),	 -- 542	7
	 ("00000000000000000000000000000110"),	 -- 541	6
	 ("00000000000000000000000000000101"),	 -- 540	5
	 ("00000000000000000000000000000100"),	 -- 539	4
	 ("00000000000000000000000000000011"),	 -- 538	3
	 ("00000000000000000000000000000010"),	 -- 537	2
	 ("00000000000000000000000000000001"),	 -- 536	1
	 ("00000000000000000000000000001000"),	 -- 535	8
	 ("00000000000000000000000000000111"),	 -- 534	7
	 ("00000000000000000000000000000110"),	 -- 533	6
	 ("00000000000000000000000000000101"),	 -- 532	5
	 ("00000000000000000000000000000100"),	 -- 531	4
	 ("00000000000000000000000000000011"),	 -- 530	3
	 ("00000000000000000000000000000010"),	 -- 529	2
	 ("00000000000000000000000000000001"),	 -- 528	1
	 ("00000000000000000000000000001000"),	 -- 527	8
	 ("00000000000000000000000000000111"),	 -- 526	7
	 ("00000000000000000000000000000110"),	 -- 525	6
	 ("00000000000000000000000000000101"),	 -- 524	5
	 ("00000000000000000000000000000100"),	 -- 523	4
	 ("00000000000000000000000000000011"),	 -- 522	3
	 ("00000000000000000000000000000010"),	 -- 521	2
	 ("00000000000000000000000000000001"),	 -- 520	1
	 ("00000000000000000000000000001000"),	 -- 519	8
	 ("00000000000000000000000000000111"),	 -- 518	7
	 ("00000000000000000000000000000110"),	 -- 517	6
	 ("00000000000000000000000000000101"),	 -- 516	5
	 ("00000000000000000000000000000100"),	 -- 515	4
	 ("00000000000000000000000000000011"),	 -- 514	3
	 ("00000000000000000000000000000010"),	 -- 513	2
	 ("00000000000000000000000000000001"),	 -- 512	1
	 ("00000000000000000000000000001000"),	 -- 511	8
	 ("00000000000000000000000000000111"),	 -- 510	7
	 ("00000000000000000000000000000110"),	 -- 509	6
	 ("00000000000000000000000000000101"),	 -- 508	5
	 ("00000000000000000000000000000100"),	 -- 507	4
	 ("00000000000000000000000000000011"),	 -- 506	3
	 ("00000000000000000000000000000010"),	 -- 505	2
	 ("00000000000000000000000000000001"),	 -- 504	1
	 ("00000000000000000000000000001000"),	 -- 503	8
	 ("00000000000000000000000000000111"),	 -- 502	7
	 ("00000000000000000000000000000110"),	 -- 501	6
	 ("00000000000000000000000000000101"),	 -- 500	5
	 ("00000000000000000000000000000100"),	 -- 499	4
	 ("00000000000000000000000000000011"),	 -- 498	3
	 ("00000000000000000000000000000010"),	 -- 497	2
	 ("00000000000000000000000000000001"),	 -- 496	1
	 ("00000000000000000000000000001000"),	 -- 495	8
	 ("00000000000000000000000000000111"),	 -- 494	7
	 ("00000000000000000000000000000110"),	 -- 493	6
	 ("00000000000000000000000000000101"),	 -- 492	5
	 ("00000000000000000000000000000100"),	 -- 491	4
	 ("00000000000000000000000000000011"),	 -- 490	3
	 ("00000000000000000000000000000010"),	 -- 489	2
	 ("00000000000000000000000000000001"),	 -- 488	1
	 ("00000000000000000000000000001000"),	 -- 487	8
	 ("00000000000000000000000000000111"),	 -- 486	7
	 ("00000000000000000000000000000110"),	 -- 485	6
	 ("00000000000000000000000000000101"),	 -- 484	5
	 ("00000000000000000000000000000100"),	 -- 483	4
	 ("00000000000000000000000000000011"),	 -- 482	3
	 ("00000000000000000000000000000010"),	 -- 481	2
	 ("00000000000000000000000000000001"),	 -- 480	1
	 ("00000000000000000000000000001000"),	 -- 479	8
	 ("00000000000000000000000000000111"),	 -- 478	7
	 ("00000000000000000000000000000110"),	 -- 477	6
	 ("00000000000000000000000000000101"),	 -- 476	5
	 ("00000000000000000000000000000100"),	 -- 475	4
	 ("00000000000000000000000000000011"),	 -- 474	3
	 ("00000000000000000000000000000010"),	 -- 473	2
	 ("00000000000000000000000000000001"),	 -- 472	1
	 ("00000000000000000000000000001000"),	 -- 471	8
	 ("00000000000000000000000000000111"),	 -- 470	7
	 ("00000000000000000000000000000110"),	 -- 469	6
	 ("00000000000000000000000000000101"),	 -- 468	5
	 ("00000000000000000000000000000100"),	 -- 467	4
	 ("00000000000000000000000000000011"),	 -- 466	3
	 ("00000000000000000000000000000010"),	 -- 465	2
	 ("00000000000000000000000000000001"),	 -- 464	1
	 ("00000000000000000000000000001000"),	 -- 463	8
	 ("00000000000000000000000000000111"),	 -- 462	7
	 ("00000000000000000000000000000110"),	 -- 461	6
	 ("00000000000000000000000000000101"),	 -- 460	5
	 ("00000000000000000000000000000100"),	 -- 459	4
	 ("00000000000000000000000000000011"),	 -- 458	3
	 ("00000000000000000000000000000010"),	 -- 457	2
	 ("00000000000000000000000000000001"),	 -- 456	1
	 ("00000000000000000000000000001000"),	 -- 455	8
	 ("00000000000000000000000000000111"),	 -- 454	7
	 ("00000000000000000000000000000110"),	 -- 453	6
	 ("00000000000000000000000000000101"),	 -- 452	5
	 ("00000000000000000000000000000100"),	 -- 451	4
	 ("00000000000000000000000000000011"),	 -- 450	3
	 ("00000000000000000000000000000010"),	 -- 449	2
	 ("00000000000000000000000000000001"),	 -- 448	1
	 ("00000000000000000000000000001000"),	 -- 447	8
	 ("00000000000000000000000000000111"),	 -- 446	7
	 ("00000000000000000000000000000110"),	 -- 445	6
	 ("00000000000000000000000000000101"),	 -- 444	5
	 ("00000000000000000000000000000100"),	 -- 443	4
	 ("00000000000000000000000000000011"),	 -- 442	3
	 ("00000000000000000000000000000010"),	 -- 441	2
	 ("00000000000000000000000000000001"),	 -- 440	1
	 ("00000000000000000000000000001000"),	 -- 439	8
	 ("00000000000000000000000000000111"),	 -- 438	7
	 ("00000000000000000000000000000110"),	 -- 437	6
	 ("00000000000000000000000000000101"),	 -- 436	5
	 ("00000000000000000000000000000100"),	 -- 435	4
	 ("00000000000000000000000000000011"),	 -- 434	3
	 ("00000000000000000000000000000010"),	 -- 433	2
	 ("00000000000000000000000000000001"),	 -- 432	1
	 ("00000000000000000000000000001000"),	 -- 431	8
	 ("00000000000000000000000000000111"),	 -- 430	7
	 ("00000000000000000000000000000110"),	 -- 429	6
	 ("00000000000000000000000000000101"),	 -- 428	5
	 ("00000000000000000000000000000100"),	 -- 427	4
	 ("00000000000000000000000000000011"),	 -- 426	3
	 ("00000000000000000000000000000010"),	 -- 425	2
	 ("00000000000000000000000000000001"),	 -- 424	1
	 ("00000000000000000000000000001000"),	 -- 423	8
	 ("00000000000000000000000000000111"),	 -- 422	7
	 ("00000000000000000000000000000110"),	 -- 421	6
	 ("00000000000000000000000000000101"),	 -- 420	5
	 ("00000000000000000000000000000100"),	 -- 419	4
	 ("00000000000000000000000000000011"),	 -- 418	3
	 ("00000000000000000000000000000010"),	 -- 417	2
	 ("00000000000000000000000000000001"),	 -- 416	1
	 ("00000000000000000000000000001000"),	 -- 415	8
	 ("00000000000000000000000000000111"),	 -- 414	7
	 ("00000000000000000000000000000110"),	 -- 413	6
	 ("00000000000000000000000000000101"),	 -- 412	5
	 ("00000000000000000000000000000100"),	 -- 411	4
	 ("00000000000000000000000000000011"),	 -- 410	3
	 ("00000000000000000000000000000010"),	 -- 409	2
	 ("00000000000000000000000000000001"),	 -- 408	1
	 ("00000000000000000000000000001000"),	 -- 407	8
	 ("00000000000000000000000000000111"),	 -- 406	7
	 ("00000000000000000000000000000110"),	 -- 405	6
	 ("00000000000000000000000000000101"),	 -- 404	5
	 ("00000000000000000000000000000100"),	 -- 403	4
	 ("00000000000000000000000000000011"),	 -- 402	3
	 ("00000000000000000000000000000010"),	 -- 401	2
	 ("00000000000000000000000000000001"),	 -- 400	1
	 ("00000000000000000000000000001000"),	 -- 399	8
	 ("00000000000000000000000000000111"),	 -- 398	7
	 ("00000000000000000000000000000110"),	 -- 397	6
	 ("00000000000000000000000000000101"),	 -- 396	5
	 ("00000000000000000000000000000100"),	 -- 395	4
	 ("00000000000000000000000000000011"),	 -- 394	3
	 ("00000000000000000000000000000010"),	 -- 393	2
	 ("00000000000000000000000000000001"),	 -- 392	1
	 ("00000000000000000000000000001000"),	 -- 391	8
	 ("00000000000000000000000000000111"),	 -- 390	7
	 ("00000000000000000000000000000110"),	 -- 389	6
	 ("00000000000000000000000000000101"),	 -- 388	5
	 ("00000000000000000000000000000100"),	 -- 387	4
	 ("00000000000000000000000000000011"),	 -- 386	3
	 ("00000000000000000000000000000010"),	 -- 385	2
	 ("00000000000000000000000000000001"),	 -- 384	1
	 ("00000000000000000000000000001000"),	 -- 383	8
	 ("00000000000000000000000000000111"),	 -- 382	7
	 ("00000000000000000000000000000110"),	 -- 381	6
	 ("00000000000000000000000000000101"),	 -- 380	5
	 ("00000000000000000000000000000100"),	 -- 379	4
	 ("00000000000000000000000000000011"),	 -- 378	3
	 ("00000000000000000000000000000010"),	 -- 377	2
	 ("00000000000000000000000000000001"),	 -- 376	1
	 ("00000000000000000000000000001000"),	 -- 375	8
	 ("00000000000000000000000000000111"),	 -- 374	7
	 ("00000000000000000000000000000110"),	 -- 373	6
	 ("00000000000000000000000000000101"),	 -- 372	5
	 ("00000000000000000000000000000100"),	 -- 371	4
	 ("00000000000000000000000000000011"),	 -- 370	3
	 ("00000000000000000000000000000010"),	 -- 369	2
	 ("00000000000000000000000000000001"),	 -- 368	1
	 ("00000000000000000000000000001000"),	 -- 367	8
	 ("00000000000000000000000000000111"),	 -- 366	7
	 ("00000000000000000000000000000110"),	 -- 365	6
	 ("00000000000000000000000000000101"),	 -- 364	5
	 ("00000000000000000000000000000100"),	 -- 363	4
	 ("00000000000000000000000000000011"),	 -- 362	3
	 ("00000000000000000000000000000010"),	 -- 361	2
	 ("00000000000000000000000000000001"),	 -- 360	1
	 ("00000000000000000000000000001000"),	 -- 359	8
	 ("00000000000000000000000000000111"),	 -- 358	7
	 ("00000000000000000000000000000110"),	 -- 357	6
	 ("00000000000000000000000000000101"),	 -- 356	5
	 ("00000000000000000000000000000100"),	 -- 355	4
	 ("00000000000000000000000000000011"),	 -- 354	3
	 ("00000000000000000000000000000010"),	 -- 353	2
	 ("00000000000000000000000000000001"),	 -- 352	1
	 ("00000000000000000000000000001000"),	 -- 351	8
	 ("00000000000000000000000000000111"),	 -- 350	7
	 ("00000000000000000000000000000110"),	 -- 349	6
	 ("00000000000000000000000000000101"),	 -- 348	5
	 ("00000000000000000000000000000100"),	 -- 347	4
	 ("00000000000000000000000000000011"),	 -- 346	3
	 ("00000000000000000000000000000010"),	 -- 345	2
	 ("00000000000000000000000000000001"),	 -- 344	1
	 ("00000000000000000000000000001000"),	 -- 343	8
	 ("00000000000000000000000000000111"),	 -- 342	7
	 ("00000000000000000000000000000110"),	 -- 341	6
	 ("00000000000000000000000000000101"),	 -- 340	5
	 ("00000000000000000000000000000100"),	 -- 339	4
	 ("00000000000000000000000000000011"),	 -- 338	3
	 ("00000000000000000000000000000010"),	 -- 337	2
	 ("00000000000000000000000000000001"),	 -- 336	1
	 ("00000000000000000000000000001000"),	 -- 335	8
	 ("00000000000000000000000000000111"),	 -- 334	7
	 ("00000000000000000000000000000110"),	 -- 333	6
	 ("00000000000000000000000000000101"),	 -- 332	5
	 ("00000000000000000000000000000100"),	 -- 331	4
	 ("00000000000000000000000000000011"),	 -- 330	3
	 ("00000000000000000000000000000010"),	 -- 329	2
	 ("00000000000000000000000000000001"),	 -- 328	1
	 ("00000000000000000000000000001000"),	 -- 327	8
	 ("00000000000000000000000000000111"),	 -- 326	7
	 ("00000000000000000000000000000110"),	 -- 325	6
	 ("00000000000000000000000000000101"),	 -- 324	5
	 ("00000000000000000000000000000100"),	 -- 323	4
	 ("00000000000000000000000000000011"),	 -- 322	3
	 ("00000000000000000000000000000010"),	 -- 321	2
	 ("00000000000000000000000000000001"),	 -- 320	1
	 ("00000000000000000000000000001000"),	 -- 319	8
	 ("00000000000000000000000000000111"),	 -- 318	7
	 ("00000000000000000000000000000110"),	 -- 317	6
	 ("00000000000000000000000000000101"),	 -- 316	5
	 ("00000000000000000000000000000100"),	 -- 315	4
	 ("00000000000000000000000000000011"),	 -- 314	3
	 ("00000000000000000000000000000010"),	 -- 313	2
	 ("00000000000000000000000000000001"),	 -- 312	1
	 ("00000000000000000000000000001000"),	 -- 311	8
	 ("00000000000000000000000000000111"),	 -- 310	7
	 ("00000000000000000000000000000110"),	 -- 309	6
	 ("00000000000000000000000000000101"),	 -- 308	5
	 ("00000000000000000000000000000100"),	 -- 307	4
	 ("00000000000000000000000000000011"),	 -- 306	3
	 ("00000000000000000000000000000010"),	 -- 305	2
	 ("00000000000000000000000000000001"),	 -- 304	1
	 ("00000000000000000000000000001000"),	 -- 303	8
	 ("00000000000000000000000000000111"),	 -- 302	7
	 ("00000000000000000000000000000110"),	 -- 301	6
	 ("00000000000000000000000000000101"),	 -- 300	5
	 ("00000000000000000000000000000100"),	 -- 299	4
	 ("00000000000000000000000000000011"),	 -- 298	3
	 ("00000000000000000000000000000010"),	 -- 297	2
	 ("00000000000000000000000000000001"),	 -- 296	1
	 ("00000000000000000000000000001000"),	 -- 295	8
	 ("00000000000000000000000000000111"),	 -- 294	7
	 ("00000000000000000000000000000110"),	 -- 293	6
	 ("00000000000000000000000000000101"),	 -- 292	5
	 ("00000000000000000000000000000100"),	 -- 291	4
	 ("00000000000000000000000000000011"),	 -- 290	3
	 ("00000000000000000000000000000010"),	 -- 289	2
	 ("00000000000000000000000000000001"),	 -- 288	1
	 ("00000000000000000000000000001000"),	 -- 287	8
	 ("00000000000000000000000000000111"),	 -- 286	7
	 ("00000000000000000000000000000110"),	 -- 285	6
	 ("00000000000000000000000000000101"),	 -- 284	5
	 ("00000000000000000000000000000100"),	 -- 283	4
	 ("00000000000000000000000000000011"),	 -- 282	3
	 ("00000000000000000000000000000010"),	 -- 281	2
	 ("00000000000000000000000000000001"),	 -- 280	1
	 ("00000000000000000000000000001000"),	 -- 279	8
	 ("00000000000000000000000000000111"),	 -- 278	7
	 ("00000000000000000000000000000110"),	 -- 277	6
	 ("00000000000000000000000000000101"),	 -- 276	5
	 ("00000000000000000000000000000100"),	 -- 275	4
	 ("00000000000000000000000000000011"),	 -- 274	3
	 ("00000000000000000000000000000010"),	 -- 273	2
	 ("00000000000000000000000000000001"),	 -- 272	1
	 ("00000000000000000000000000001000"),	 -- 271	8
	 ("00000000000000000000000000000111"),	 -- 270	7
	 ("00000000000000000000000000000110"),	 -- 269	6
	 ("00000000000000000000000000000101"),	 -- 268	5
	 ("00000000000000000000000000000100"),	 -- 267	4
	 ("00000000000000000000000000000011"),	 -- 266	3
	 ("00000000000000000000000000000010"),	 -- 265	2
	 ("00000000000000000000000000000001"),	 -- 264	1
	 ("00000000000000000000000000001000"),	 -- 263	8
	 ("00000000000000000000000000000111"),	 -- 262	7
	 ("00000000000000000000000000000110"),	 -- 261	6
	 ("00000000000000000000000000000101"),	 -- 260	5
	 ("00000000000000000000000000000100"),	 -- 259	4
	 ("00000000000000000000000000000011"),	 -- 258	3
	 ("00000000000000000000000000000010"),	 -- 257	2
	 ("00000000000000000000000000000001"),	 -- 256	1
	 ("00000000000000000000000000001000"),	 -- 255	8
	 ("00000000000000000000000000000111"),	 -- 254	7
	 ("00000000000000000000000000000110"),	 -- 253	6
	 ("00000000000000000000000000000101"),	 -- 252	5
	 ("00000000000000000000000000000100"),	 -- 251	4
	 ("00000000000000000000000000000011"),	 -- 250	3
	 ("00000000000000000000000000000010"),	 -- 249	2
	 ("00000000000000000000000000000001"),	 -- 248	1
	 ("00000000000000000000000000001000"),	 -- 247	8
	 ("00000000000000000000000000000111"),	 -- 246	7
	 ("00000000000000000000000000000110"),	 -- 245	6
	 ("00000000000000000000000000000101"),	 -- 244	5
	 ("00000000000000000000000000000100"),	 -- 243	4
	 ("00000000000000000000000000000011"),	 -- 242	3
	 ("00000000000000000000000000000010"),	 -- 241	2
	 ("00000000000000000000000000000001"),	 -- 240	1
	 ("00000000000000000000000000001000"),	 -- 239	8
	 ("00000000000000000000000000000111"),	 -- 238	7
	 ("00000000000000000000000000000110"),	 -- 237	6
	 ("00000000000000000000000000000101"),	 -- 236	5
	 ("00000000000000000000000000000100"),	 -- 235	4
	 ("00000000000000000000000000000011"),	 -- 234	3
	 ("00000000000000000000000000000010"),	 -- 233	2
	 ("00000000000000000000000000000001"),	 -- 232	1
	 ("00000000000000000000000000001000"),	 -- 231	8
	 ("00000000000000000000000000000111"),	 -- 230	7
	 ("00000000000000000000000000000110"),	 -- 229	6
	 ("00000000000000000000000000000101"),	 -- 228	5
	 ("00000000000000000000000000000100"),	 -- 227	4
	 ("00000000000000000000000000000011"),	 -- 226	3
	 ("00000000000000000000000000000010"),	 -- 225	2
	 ("00000000000000000000000000000001"),	 -- 224	1
	 ("00000000000000000000000000001000"),	 -- 223	8
	 ("00000000000000000000000000000111"),	 -- 222	7
	 ("00000000000000000000000000000110"),	 -- 221	6
	 ("00000000000000000000000000000101"),	 -- 220	5
	 ("00000000000000000000000000000100"),	 -- 219	4
	 ("00000000000000000000000000000011"),	 -- 218	3
	 ("00000000000000000000000000000010"),	 -- 217	2
	 ("00000000000000000000000000000001"),	 -- 216	1
	 ("00000000000000000000000000001000"),	 -- 215	8
	 ("00000000000000000000000000000111"),	 -- 214	7
	 ("00000000000000000000000000000110"),	 -- 213	6
	 ("00000000000000000000000000000101"),	 -- 212	5
	 ("00000000000000000000000000000100"),	 -- 211	4
	 ("00000000000000000000000000000011"),	 -- 210	3
	 ("00000000000000000000000000000010"),	 -- 209	2
	 ("00000000000000000000000000000001"),	 -- 208	1
	 ("00000000000000000000000000001000"),	 -- 207	8
	 ("00000000000000000000000000000111"),	 -- 206	7
	 ("00000000000000000000000000000110"),	 -- 205	6
	 ("00000000000000000000000000000101"),	 -- 204	5
	 ("00000000000000000000000000000100"),	 -- 203	4
	 ("00000000000000000000000000000011"),	 -- 202	3
	 ("00000000000000000000000000000010"),	 -- 201	2
	 ("00000000000000000000000000000001"),	 -- 200	1
	 ("00000000000000000000000000001000"),	 -- 199	8
	 ("00000000000000000000000000000111"),	 -- 198	7
	 ("00000000000000000000000000000110"),	 -- 197	6
	 ("00000000000000000000000000000101"),	 -- 196	5
	 ("00000000000000000000000000000100"),	 -- 195	4
	 ("00000000000000000000000000000011"),	 -- 194	3
	 ("00000000000000000000000000000010"),	 -- 193	2
	 ("00000000000000000000000000000001"),	 -- 192	1
	 ("00000000000000000000000000001000"),	 -- 191	8
	 ("00000000000000000000000000000111"),	 -- 190	7
	 ("00000000000000000000000000000110"),	 -- 189	6
	 ("00000000000000000000000000000101"),	 -- 188	5
	 ("00000000000000000000000000000100"),	 -- 187	4
	 ("00000000000000000000000000000011"),	 -- 186	3
	 ("00000000000000000000000000000010"),	 -- 185	2
	 ("00000000000000000000000000000001"),	 -- 184	1
	 ("00000000000000000000000000001000"),	 -- 183	8
	 ("00000000000000000000000000000111"),	 -- 182	7
	 ("00000000000000000000000000000110"),	 -- 181	6
	 ("00000000000000000000000000000101"),	 -- 180	5
	 ("00000000000000000000000000000100"),	 -- 179	4
	 ("00000000000000000000000000000011"),	 -- 178	3
	 ("00000000000000000000000000000010"),	 -- 177	2
	 ("00000000000000000000000000000001"),	 -- 176	1
	 ("00000000000000000000000000001000"),	 -- 175	8
	 ("00000000000000000000000000000111"),	 -- 174	7
	 ("00000000000000000000000000000110"),	 -- 173	6
	 ("00000000000000000000000000000101"),	 -- 172	5
	 ("00000000000000000000000000000100"),	 -- 171	4
	 ("00000000000000000000000000000011"),	 -- 170	3
	 ("00000000000000000000000000000010"),	 -- 169	2
	 ("00000000000000000000000000000001"),	 -- 168	1
	 ("00000000000000000000000000001000"),	 -- 167	8
	 ("00000000000000000000000000000111"),	 -- 166	7
	 ("00000000000000000000000000000110"),	 -- 165	6
	 ("00000000000000000000000000000101"),	 -- 164	5
	 ("00000000000000000000000000000100"),	 -- 163	4
	 ("00000000000000000000000000000011"),	 -- 162	3
	 ("00000000000000000000000000000010"),	 -- 161	2
	 ("00000000000000000000000000000001"),	 -- 160	1
	 ("00000000000000000000000000001000"),	 -- 159	8
	 ("00000000000000000000000000000111"),	 -- 158	7
	 ("00000000000000000000000000000110"),	 -- 157	6
	 ("00000000000000000000000000000101"),	 -- 156	5
	 ("00000000000000000000000000000100"),	 -- 155	4
	 ("00000000000000000000000000000011"),	 -- 154	3
	 ("00000000000000000000000000000010"),	 -- 153	2
	 ("00000000000000000000000000000001"),	 -- 152	1
	 ("00000000000000000000000000001000"),	 -- 151	8
	 ("00000000000000000000000000000111"),	 -- 150	7
	 ("00000000000000000000000000000110"),	 -- 149	6
	 ("00000000000000000000000000000101"),	 -- 148	5
	 ("00000000000000000000000000000100"),	 -- 147	4
	 ("00000000000000000000000000000011"),	 -- 146	3
	 ("00000000000000000000000000000010"),	 -- 145	2
	 ("00000000000000000000000000000001"),	 -- 144	1
	 ("00000000000000000000000000001000"),	 -- 143	8
	 ("00000000000000000000000000000111"),	 -- 142	7
	 ("00000000000000000000000000000110"),	 -- 141	6
	 ("00000000000000000000000000000101"),	 -- 140	5
	 ("00000000000000000000000000000100"),	 -- 139	4
	 ("00000000000000000000000000000011"),	 -- 138	3
	 ("00000000000000000000000000000010"),	 -- 137	2
	 ("00000000000000000000000000000001"),	 -- 136	1
	 ("00000000000000000000000000001000"),	 -- 135	8
	 ("00000000000000000000000000000111"),	 -- 134	7
	 ("00000000000000000000000000000110"),	 -- 133	6
	 ("00000000000000000000000000000101"),	 -- 132	5
	 ("00000000000000000000000000000100"),	 -- 131	4
	 ("00000000000000000000000000000011"),	 -- 130	3
	 ("00000000000000000000000000000010"),	 -- 129	2
	 ("00000000000000000000000000000001"),	 -- 128	1
	 ("00000000000000000000000000001000"),	 -- 127	8
	 ("00000000000000000000000000000111"),	 -- 126	7
	 ("00000000000000000000000000000110"),	 -- 125	6
	 ("00000000000000000000000000000101"),	 -- 124	5
	 ("00000000000000000000000000000100"),	 -- 123	4
	 ("00000000000000000000000000000011"),	 -- 122	3
	 ("00000000000000000000000000000010"),	 -- 121	2
	 ("00000000000000000000000000000001"),	 -- 120	1
	 ("00000000000000000000000000001000"),	 -- 119	8
	 ("00000000000000000000000000000111"),	 -- 118	7
	 ("00000000000000000000000000000110"),	 -- 117	6
	 ("00000000000000000000000000000101"),	 -- 116	5
	 ("00000000000000000000000000000100"),	 -- 115	4
	 ("00000000000000000000000000000011"),	 -- 114	3
	 ("00000000000000000000000000000010"),	 -- 113	2
	 ("00000000000000000000000000000001"),	 -- 112	1
	 ("00000000000000000000000000001000"),	 -- 111	8
	 ("00000000000000000000000000000111"),	 -- 110	7
	 ("00000000000000000000000000000110"),	 -- 109	6
	 ("00000000000000000000000000000101"),	 -- 108	5
	 ("00000000000000000000000000000100"),	 -- 107	4
	 ("00000000000000000000000000000011"),	 -- 106	3
	 ("00000000000000000000000000000010"),	 -- 105	2
	 ("00000000000000000000000000000001"),	 -- 104	1
	 ("00000000000000000000000000001000"),	 -- 103	8
	 ("00000000000000000000000000000111"),	 -- 102	7
	 ("00000000000000000000000000000110"),	 -- 101	6
	 ("00000000000000000000000000000101"),	 -- 100	5
	 ("00000000000000000000000000000100"),	 -- 99	4
	 ("00000000000000000000000000000011"),	 -- 98	3
	 ("00000000000000000000000000000010"),	 -- 97	2
	 ("00000000000000000000000000000001"),	 -- 96	1
	 ("00000000000000000000000000001000"),	 -- 95	8
	 ("00000000000000000000000000000111"),	 -- 94	7
	 ("00000000000000000000000000000110"),	 -- 93	6
	 ("00000000000000000000000000000101"),	 -- 92	5
	 ("00000000000000000000000000000100"),	 -- 91	4
	 ("00000000000000000000000000000011"),	 -- 90	3
	 ("00000000000000000000000000000010"),	 -- 89	2
	 ("00000000000000000000000000000001"),	 -- 88	1
	 ("00000000000000000000000000001000"),	 -- 87	8
	 ("00000000000000000000000000000111"),	 -- 86	7
	 ("00000000000000000000000000000110"),	 -- 85	6
	 ("00000000000000000000000000000101"),	 -- 84	5
	 ("00000000000000000000000000000100"),	 -- 83	4
	 ("00000000000000000000000000000011"),	 -- 82	3
	 ("00000000000000000000000000000010"),	 -- 81	2
	 ("00000000000000000000000000000001"),	 -- 80	1
	 ("00000000000000000000000000001000"),	 -- 79	8
	 ("00000000000000000000000000000111"),	 -- 78	7
	 ("00000000000000000000000000000110"),	 -- 77	6
	 ("00000000000000000000000000000101"),	 -- 76	5
	 ("00000000000000000000000000000100"),	 -- 75	4
	 ("00000000000000000000000000000011"),	 -- 74	3
	 ("00000000000000000000000000000010"),	 -- 73	2
	 ("00000000000000000000000000000001"),	 -- 72	1
	 ("00000000000000000000000000001000"),	 -- 71	8
	 ("00000000000000000000000000000111"),	 -- 70	7
	 ("00000000000000000000000000000110"),	 -- 69	6
	 ("00000000000000000000000000000101"),	 -- 68	5
	 ("00000000000000000000000000000100"),	 -- 67	4
	 ("00000000000000000000000000000011"),	 -- 66	3
	 ("00000000000000000000000000000010"),	 -- 65	2
	 ("00000000000000000000000000000001"),	 -- 64	1
	 ("00000000000000000000000000001000"),	 -- 63	8
	 ("00000000000000000000000000000111"),	 -- 62	7
	 ("00000000000000000000000000000110"),	 -- 61	6
	 ("00000000000000000000000000000101"),	 -- 60	5
	 ("00000000000000000000000000000100"),	 -- 59	4
	 ("00000000000000000000000000000011"),	 -- 58	3
	 ("00000000000000000000000000000010"),	 -- 57	2
	 ("00000000000000000000000000000001"),	 -- 56	1
	 ("00000000000000000000000000001000"),	 -- 55	8
	 ("00000000000000000000000000000111"),	 -- 54	7
	 ("00000000000000000000000000000110"),	 -- 53	6
	 ("00000000000000000000000000000101"),	 -- 52	5
	 ("00000000000000000000000000000100"),	 -- 51	4
	 ("00000000000000000000000000000011"),	 -- 50	3
	 ("00000000000000000000000000000010"),	 -- 49	2
	 ("00000000000000000000000000000001"),	 -- 48	1
	 ("00000000000000000000000000001000"),	 -- 47	8
	 ("00000000000000000000000000000111"),	 -- 46	7
	 ("00000000000000000000000000000110"),	 -- 45	6
	 ("00000000000000000000000000000101"),	 -- 44	5
	 ("00000000000000000000000000000100"),	 -- 43	4
	 ("00000000000000000000000000000011"),	 -- 42	3
	 ("00000000000000000000000000000010"),	 -- 41	2
	 ("00000000000000000000000000000001"),	 -- 40	1
	 ("00000000000000000000000000001000"),	 -- 39	8
	 ("00000000000000000000000000000111"),	 -- 38	7
	 ("00000000000000000000000000000110"),	 -- 37	6
	 ("00000000000000000000000000000101"),	 -- 36	5
	 ("00000000000000000000000000000100"),	 -- 35	4
	 ("00000000000000000000000000000011"),	 -- 34	3
	 ("00000000000000000000000000000010"),	 -- 33	2
	 ("00000000000000000000000000000001"),	 -- 32	1
	 ("00000000000000000000000000001000"),	 -- 31	8
	 ("00000000000000000000000000000111"),	 -- 30	7
	 ("00000000000000000000000000000110"),	 -- 29	6
	 ("00000000000000000000000000000101"),	 -- 28	5
	 ("00000000000000000000000000000100"),	 -- 27	4
	 ("00000000000000000000000000000011"),	 -- 26	3
	 ("00000000000000000000000000000010"),	 -- 25	2
	 ("00000000000000000000000000000001"),	 -- 24	1
	 ("00000000000000000000000000001000"),	 -- 23	8
	 ("00000000000000000000000000000111"),	 -- 22	7
	 ("00000000000000000000000000000110"),	 -- 21	6
	 ("00000000000000000000000000000101"),	 -- 20	5
	 ("00000000000000000000000000000100"),	 -- 19	4
	 ("00000000000000000000000000000011"),	 -- 18	3
	 ("00000000000000000000000000000010"),	 -- 17	2
	 ("00000000000000000000000000000001"),	 -- 16	1
	 ("00000000000000000000000000001000"),	 -- 15	8
	 ("00000000000000000000000000000111"),	 -- 14	7
	 ("00000000000000000000000000000110"),	 -- 13	6
	 ("00000000000000000000000000000101"),	 -- 12	5
	 ("00000000000000000000000000000100"),	 -- 11	4
	 ("00000000000000000000000000000011"),	 -- 10	3
	 ("00000000000000000000000000000010"),	 -- 9	2
	 ("00000000000000000000000000000001"),	 -- 8	1
	 ("00000000000000000000000000001000"),	 -- 7	8
	 ("00000000000000000000000000000111"),	 -- 6	7
	 ("00000000000000000000000000000110"),	 -- 5	6
	 ("00000000000000000000000000000101"),	 -- 4	5
	 ("00000000000000000000000000000100"),	 -- 3	4
	 ("00000000000000000000000000000011"),	 -- 2	3
	 ("00000000000000000000000000000010"),	 -- 1	2
	 ("00000000000000000000000000000001"));	 -- 0	1

begin
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we = '1') then
        RAM(conv_integer(address)) <= data_in;
        data_out <= RAM(conv_integer(read_a));
      elsif (oe = '1') then
        data_out <= RAM(conv_integer(read_a));
      end if;
      read_a <= address;
    end if;
  end process;
end rtl;
